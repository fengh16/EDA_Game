// clk为控制的时钟信号，周期性输出0和1。在这里给一个输入信号，让这个module工作。
module generator_1000hz(c, clk);
	input c;
	output reg clk;
	reg [31:0] cnt;
	parameter period = 40000;

	initial
		clk = 0;
	
	always @ (posedge c) begin
		if (cnt == (period >> 1) - 1) begin
			clk <= 1'b1;
			cnt <= cnt + 1;
		end else if (cnt == period - 1) begin
			clk <= 1'b0;
			cnt <= 0;
		end else
			cnt <= cnt + 1;
	end
endmodule

// 每次时钟切换，就换不同的数码管显示。因为频率很高，就不会让人发现闪烁。
module counter_scan(clk, scan_cnt);
	input clk;
	output reg [2:0] scan_cnt;

	initial
		scan_cnt <= 0;

	always @(posedge clk) begin
		if (scan_cnt == 3'd5)
			scan_cnt <= 3'd0;
		else
			scan_cnt <= scan_cnt + 3'd1;
	end
endmodule

// 选择数码管显示的时候，将刚才上面那个函数的输出换到数码管选通的控制
module selector_digit(scan_cnt, digit);
	input [2:0] scan_cnt;
	output reg [1:6] digit;
	
	always @ (scan_cnt)
		case (scan_cnt)
			0: digit <= 6'b111110;
			1: digit <= 6'b111101;
			2: digit <= 6'b111011;
			3: digit <= 6'b110111;
			4: digit <= 6'b101111;
			5: digit <= 6'b011111;
			default: digit <= 6'b111111;
		endcase
endmodule

// 把所有数码管应该输出的东西放在这里，然后就可以通过scan_cnt来控制哪个要输出
module selector_seg(scan_cnt, dig1, dig2, dig3, dig4, dig5, dig6, seg);
	input [2:0] scan_cnt;
	input [6:0] dig1, dig2, dig3, dig4, dig5, dig6;
	output reg [6:0] seg;
	
	always @ (scan_cnt, dig1, dig2, dig3, dig4, dig5, dig6) begin 
		case (scan_cnt)
			0: seg <= dig1;
			1: seg <= dig2;
			2: seg <= dig3;
			3: seg <= dig4;
			4: seg <= dig5;
			5: seg <= dig6;
		endcase
	end
endmodule

module Game(c, start, button, switch, speed, L, SEGNum, LED);
	input c;
	input start;
	input [2:0]button;
	input [5:0]switch;
	input [1:0]speed;
	output reg [7:0]LED;
	output [6:0]L; // Hex light output(one bit hex number);
	output [5:0]SEGNum; // Use it to determine which to light;
	wire [2:0]scan_cnt;
	wire clk;

	reg [16383:0]data1;
	reg [16383:0]data2;
	reg [16383:0]data3;

	reg [14:0]num;
	reg started;
	reg startlast;
	reg [11:0]score;

	reg [6:0]show5;
	reg [6:0]show4;
	reg [6:0]show3;
	reg [6:0]show2;
	reg [6:0]show1;
	reg [6:0]show0;

	reg [10:0]state;
	reg left;
	reg middle;
	reg right;
	reg [3:0]out;
	 
	 reg button0Last;
	 reg button1Last;
	 reg button2Last;
	 
	 reg failed;

	initial
	begin
		data1[16383:0] = 16384'b0000000000000000000000010000000000000010000100000000000001000001000000000001000000000000000000001000000000000000000000100000010000000000001000000000010000000000010010000100000001000001000010101000000000000000000000000001110000000101000000000000000011000000000100000001000000100000000000010000000000000000000000000001000000000000000000000010000000000100000000000000000100000100000100000100000001000000010000000010100100000000001010000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000000010000011000000000010001000000000100000000000000000000000000000001000000000000000110000000010001000000000000000010000001001010100100001000000000000000000000010000000100000000000100000000000000001010000100100001000000000010000000001000000000000000000000000010010000000010000000000000000000000000000000001100100000100010010000000000000100000100000000001100000000100000000100000000000000110000100000000000010001000000000100000000100100000000000000000001010000000000000001001010001000000000010000000000100000000000000000000000000000000000000000000000000000000000001000001100000001000000010000010000000000000000000000001000000000100000000000000000010000001000000100000000010000000000010001000001101000000000000000000100000000001000000000010000000000000000000000000000100010000100000000000000000000000000101010000000000000000010000000101001000000001000000000000000100000000000000000000000000000010010000000010100001000000000000000100100010010000000000000000000000110100000000000001000000000000000000000000000010000001010000000000000010000000010000000000010000001000000010100000000000100000000000000000000100000000010000010000000000000000000001000011000000000110000100000000000101000000000000011000000000000000000010000000010001100000000000000000000000000000000000000000000000010000000000000000000000001000000000010000010000000000000010000000000000000000000001000000000000000000110000001000000000000000000001000000000000000000000000000001000000010100000000000000001010000010000000000000001000011000000001000000000000000000000110000000000010010000000001010000010000001000000000000000000000100011110000000000000000000000000000000000000010000010100000100000000000001010000000100000010000001100010000000000000000000010100010100001000100000000001000000000010000000000010100000000000000001010000000000010000000000010010000000000000000000000000101000000000000010000010010000010001000000100000101000001000011000000000000000001000001010000100110000010010000000000000100001000100000001000000100000000000100000101000000000000000001101010010000000000000000000001000000001100011000001000000000000000000100000000100100010010110010000000000000100000000000000000001100001001000000000011000000000000000000000100000000010100000000000000001001000100100000001000000000010000000100000010000000000000001000000000000000010010010000101000100000010000000000001000001001001000010000000000010001000100000000100000001000000001010000000000000000000000000010000001010000101001001010000000000001001100111000000100010000000000000000000000000010000100101000000000000010000100000010010010100000000000000000000000001000010000001001001010000000000101000000000100100000001000010000000000000000010000001000011000000010000000000000010000000000000001001001000111010000100000001000100000000101000010000010000000000000000010001111001000010100000010001000000000001100000100000000010000010000001100011000000000001000001000000000000000000000000001000000000010000000010010100010010110010000001000010000000001001101000000001000001000001010000000100000000010000000000100000101000000000010111100000010000000000000100000001000010000001000000000000001000000000100000000000000001000000010000001000100000010000100000000000000001000000000000000000000000000100000000010000000000010000101000100010000000001000000000000100000000000000100110000001000010110000011000001100000100000001001000000000010010010000001001000000011000000100010000000000001000000000010000001000000100010000100010000010000100000000000000000000001000000000001010100001100010000000001000000000001000000000100010010000000000001000000000100000010100101001000100000001100000000100001010001000110000000001000100100001110000000010010000000001000100000000000101000110000101010000000000000100000000000101000000000000000001000000000000000011001000000110000000000000100000001100000100000000001101000000000010000000100000100001100010000000000011000000100010001000101110000000000000000100000000010000000000000000100000100010100101001011000000000000000001110000010001001000000000011000000100000000000110000100000000001000000000000011000000100000100000000100000100000001000001100100000010100000000000000000100000000001010000000000000000000000110100001010001000000111010010000100000010110100100001000000000100000000000010000011000000100000000001010000000000010010000000011000000010010100000000100000000000000100000100001010000000000110110000000010001000100100000000000100100000000000000010010000000100000001010000101000001010110000000010110100000000000000000000100000000000000100000000000000000000110110000000010000000010000100101010010001000000000100000000000000001111001000000100010100000110000000000001000000100000000000000000000100000010101100001000010001000000000000000000001000100001000001000100000010000001000001000100110101000000010100000110000010100000000010000000100000001000000000000000010000010110011000000011100001000000100000001010001000000000000010001000000000010000000110100000000100000000000001010110000000001000000110000000001000001001011111000000000000100000010000000000110001000000000000010000000100000110000001010000001000000010100010000000001000000100000010001001000000011000000000100000000000000011101100001000010000100001000000010000000010000000001110000010000100000010000000100000000000000110010000000000000000100000011000001000000001000000100011100100100000000100000000000010000000000100000100010010000010000001000001000000001000000000100000000000000001000000010100010000000000011000000000001100001110000000000000000000000000001000000010000010001000000100000000100000010000000100100000011010010100000010010010100100000010010110100000010100000000100000000100010000000011001001010010011000000000010000000001000000001101010000000000001000011100010000000000100000000000010000001100000100010110000000011010011000100000000000001010000000101001000100000000100000101101000010001001100001000100000001010001000001010000101000000000010010010100110000000001010010010001000100000111001010001100000000000100000110000000000001001000001000000001001110000000000000011100001110000001001001000100000010000100011010000000001011000000000000000000000011000001000000000100011011101001000100001001001010010001000001100100100101010000100000000100101010000000110011110010000010000000000001100000000110001010100000010000000011001010000001000010001010100100010000000010010100000000000000000000000000001000000000101010000100101000011000000000011000111000100001010100100000001000100100000010001100010010000000000001100001000000000010000000000000000000100000010100010000000100001001000000100010010001000011011110011000110000101110010000100101100000110000010110000001000001000010010000100011111000100000000000001000001010000100000010000100000010110101000010001100011000101010000010000011000100000000010010010000110010010000010001001011000011101000000000100010000111100101000100011000001100000100000010100000000000100011010000000001000100101000110101000100100100010101000000100000101000010000101100001100110000000100010010010100000011001010001010010000010000001011011000010100001000000000000010000100010001101000000001100000000001100100100011000000001000001011000100100000000000101001000001110100001000000000001110101000000010101100001000001110011011001100000000001100110000101000010000000100001111000001010000101000010111010001000010010000100000000000000000010000010110010000000110000010000100000101000110100000000000000001000000100100000000100010000000000010010010011000110100001001011001000000100100100001100111100000000010000001000000110001100001011110010000100011000000000010000000011000010001000010111000001010100001000010010000001000000010000000000010000000010000011010000010000011010100001000000000011001010000010000011001000100100000011000001000110001000110010110100000010001000010100100110100011101001100010100101000100110000010000000010001100000001100000001100011001001001011001010000101100000110100010010000000011111010100100000000000100101000011000000000000001100010100100000000101110010101001001000011010010110000101001000010011100011111101001110100000101000100100000010111000010110110011010000111001000000010110000010010001100000010000000000001000111101001001001000010010011001100000001000000000001010011000000100001000011000000111100000001000110010001000101111001000011001100000101000110100001000001000100000000000000000101001111100000000000000101000010000101001110010010100001110001100010011000111100000010011110000100000001000001100001001100000100000001101000010000000000101111100000000000000111100000101010010001101010000000001010010110011000100101110010000110010100001101100010110010000000100000101101111000101000000100000000000001101001101110010100000100001100000101010010000000100000011000000000000100100101100100000000010010000010000100000100010000011000000100011010011100010100000100001000101010010100000000000001010011100010100010101000000100111000000100010000000000001010000010110010000010100001011001101010110010000110110000000110100000001000100110010011001100111010000000000000001000010100000011101111000010101100100100100011010001000011001000001000100011000000100000001011100000110101010011010100110101001000110001001010100000011100000100010101001001001010010100100011000010010001010000010010000000000111110001000010001000011100000000000000000101100110010001101001010000000000111100010100110000000000010011010010000000000001000100110100000000110000101000010000000001010000111010000011010100000010110010001000000100000100001000000001111100010000110110000001000010001110001010111000110010100000110010100110100001000000000010000000000101100000101101100000000100010110000001111001010100010000100100010000000000011100010010110111000010001000001001001100100010001100110000000100100100001110001000000000010000011010001000001000100100001000011000000000110010001001010110010000000011100100000010100111110010000110000010101100001000010011100000110100001000110111011101000000100001010101000110011010011100110010101100101000010001000001000101110010101011010000001101110101100001011101000110111010100010101001000000100011100100000010001011110011000000001100000000000001000000000100011000000000010010000001101001110100010111110100000101010100000001101000010100111111001111110000000011011000110000100010010000001111011010000110010100000111011000100101101000011001001110001000101110000110001001101101001000010011001000010001110001110110000101000000110100000000010010110110010001000001101100110000010110110100001011000010111000101111000100111010000100110001011110110000000010000000110001001000100100011000000110000000011010010000000001010101001010010110111011001000011100100101000100100010010010100100100011010110010110000000000101001010100000000000100011000011110000101000010000011101011000000010000110011100001000100110110000100100011101001001100000000000101110100101010100000110101100000001010001101011010001000111110011100011110000100000000100000000000010100100100000101000001011001000011111010000110010100101110000000011110000100000010001000001100011001010011011010000100001000000110100100101000100010001100110110001001111001010010000100010011000101100000000000011000011000110010000011000011000000000011000000010101000110001000000100001000110001110000001100010001100000011000101010000011000100010001010101111101100000001100001010010001000111010011000100000011100000010101110000100010010001001000100100000100100100000000010001000010000000000000010000001000001000011000100110000000011101010001100110010001000000010010000010010110011101100001000010110000101000110000011010001011110000000101100100100001010000110000100110000000001010000110011000001010000001000101100111000101001100000010111010000010110010000011001101110110010001011011100000000011100000000011110100001000100111001100011000111001100000100011111000000101110100110001011011100101001111001001100000011101000000001000001011001001011000000000101001110011100100100011000100000010100101110110000100010010000011111011101010101010010000101000110100000010110000100000100010010100010010000111110101011010011001010100011110000101010010001000001010110011101010001000100010100101010010011100000110100000100000001100011100010010000100011110001101111000010110000100001101000001111101100001101110101001000101000100010100000001000111001010000101001000000001100000000000000101101111110101010011011010000001101011010001101000000101001000101000001111010001000000001110000000001001000001111000100111010000111100010000110100100001101000001000010011101001110111011010100010101000110110011001100100000000110100101000010001101101001010101001000000101000010101100011110000001110010100110010101110001011011010001000100000000010010110111000000001110010010101010011000111010101101001011001000101100011000000010011000010001001000110010100100101001011010010110000011100100110011010101011100001001110101001111010001100100110000110111001001010110111010010100100001001111000111100110101011001001101101010001000000100000010000100110010111010011001111001000011100000110001111100110010110000000100111110110000010110000101010000000001010101111001010000100000111101011011011110001010001110110000100000011111101100000011100000000001000001111000000101110010010011000110000000000101100101001100101000110001010000110110100110001101001010000101000100000010111110001001011010011010011001110001001101100000010000101000011011110000000101100100010101001110111010100101111101100000001000110110010010010000101001001011000100100000000010111100001011101001110000111111000000001100100100110001101111000100110101011010110000001011000100010101000000000101000000100000000000101000000111100110010110000001101100100101010001101101101000001110110100110101010100001001001100000100011100110000101111000100110010001100100110110000000101000010001101111011110001110010011000011111000100001110110000101110001001000011100000010000110011001100011001001011110001000011111001110101100001011000000111000000100100110000000100101110010101001001101101001001110010100011101110001010100010100101001000101011000101100110111111110111111110100100001101000110111001110001100011100111100101000001010110111100111101011100000011111001100011011000100001111110010000011101111010010001110010001000111111000001000000010111001100010000011110011100110110001001000100000010000110100000000010000101100110000011000000100111000011100100100100101010011001011110001011000001000011001000011011100010010111011101110000111010111111000101001011110011000011111100001010010110110010011000000001010000000000110111110100011101101111000011010011110001000000011010100111011110110011001011111111100001110001010010010100100001110100000111001000000010001011110110100011111110100111100111100000101101000001111100100000100101010100010011011000001010110101110101001001111110101011010001001100000100100001010100001010100001001101111110010100011110011111011010101100011110010000010101111000001110100000000100100011111110000101101101010000001011001011001110001000100011111100101101001100110011000101100101100000100101100001100011100100101011101011001101101001011111111000111001001000010100101000100001010000111101111111101010001001001010001100100010101001111010010011100011100100010111101100101011000011100010101001001111001110001001000010110101000000101101000011000101001000110001101110001011000001001011110011100000100100010000010010111111000011010100101100111101100111011100011010001110110100011111110100110110101101111010010000001101100011000000010110001111011001011100000011010011010000011111001000100001110100001011101001001001011011001010000001100100100001000001000001100000010000001010100100010111100110111110010100110001100100110011111010111110001001000101100011000110101000101101000101000010011000001101100001100111001011100111000010101000101111110001100001111100000011101111000110010000010000100000110101111110001001001101100100111011010111000001011010000000011000000100011110001101010010111011111101101000000100001010101100111000100110110000000010000110011011111010110000010000100001010000000110100010110101101010000000011001101100101101111101000101111100100000000011001100110011010110011101000100;
		data2[16383:0] = 16384'b0000000010000000000110100000000100000000000000010000001000000000010000100000000000000000000100000100000000001100000000000000010010010001000010000100010000010011000000000000010000010100000010000000000000010010000010000001010000000001000000000000000000001000000000000000010100000000000000010000000000000000000010000000100000000010100000000000000000000000000000100000000001000000000000000001110000000000100000100000010000000000100001000010000100000000000000000000010010000010001101000000000000001000000000000000100001001001000000000000000000000000000101000010000100100100000000000000011000001010000000100101000000000000000010000000000000000000000000000000000000000000000000010000000001000000010001001000000000000000101000101000000100000000000100011001000000000000100000000000010000010000110000100000000001000000000000000000000100000010000100011000000000000000000000000010010000000001000000000000000000100100000000000000000000000000000000000100011000000000000001000000010000000000001000000001000000000000000000000001100000000000000000100000100000000000010000001001111000000000000100000000010000000000000000100000000010100000000000000010100100000000010000000000000000000000100000000000000000000000111001000000000000000000000000100000000000000000000000000010000100000000000100000000010000000000000000000000100000100000100000010000000000100000000010000000000000000000000000000010000000000000000000000100000000000010000000000010001000000000010000000000000000001000000001010000000000000000000010100010000000000000000000000000000000000000000000000000010000000110100000000000000001000000001000100000010000000000000010000100000010000000000100000100000000110000100000000100000000000010100001000000000000100000010000000000100000011000000010001000000000000000000000000000000000000100000000000000010001000000001000000000010000001001000000000100000000000000000100000010000000000000010100000000000000100000100010000010100000000000000000110000010010000000000000100000010000000100000000010000000000000000000110000010100001000000000100000000001000000000000000000000000000110000000000000000000000101000000000000000010100000011000000000000010010000001000100110000000000000000100010000010000000000000000100000000010000000000001001000000110100000000001000000000010000000010000000100110000000000010000110000000000000000000000000000001000000000000000000000000000011010000000100100010000000010011000101000000000100010010000000000100001001100011010000001100001100000010000001000000010000010000000000100000000000010000010100001000001000000010010000100000000000000001001000001000000000100000000000111000000000000001001000000001000000001000000010010000000000000100000000000110000100000000000000010110000000001000010000000000000100100110111000000000000000010000000000000010010001001011000000100000010101100000000001100000000000000000011100000001010000100000000000000001000000110010000000010000100000010000100000010100000001100000000000010000001001000100000000001000110001001010000010000000000000100000000000011100000001000010000100100010000100000001011001010000011000000100110100000101010010010100101010000000000000000000000000010100000010000000000001000000000100000110110000000100010010011000000000000101000100000000010000011000000000010000000000010001001000000000000011000110000000000000000000000000011010001001000000000100000000100000000000000000101000100000000010010000000000000000001000001000000001100000000000001010000000000000010000000001101000000011000000101110100000000000001000000000000010000000000001010000000000000010010001010000000000000000001000000011000000000000000000000100000000000000000010010000001100010000001100000001001000000100000110000000000000010000000110000000000000100000010011000010000001000000101000000000000001000000000000000000000000011010000000000010000000000000000011100000010000000000100100010100010100000100000000001000001000001000000100000001010001000100000000000000010000100000010001000000000000000001010000011000100010000000100010000000000000000000110001000001000000000001000011100010000001000100000101000000100000000000000000000000000000010000000001000010000010000000000000000000000000010010100001000000000000000100000010000000000000110000000101000000011001100100000000110000000000000000000100000000000001010100000100000011110101010000000001000000000101010001100000000100000000000000100000000000000000000000001010000000000010010010101000000001000100000010001100000000000010100100000001100000000000001000001000000000000010100011011000001000001010001001001100010000100000000100000101010000001001000000001000000000001000100000010001000000001000000000101000100001100010011001000001001000000100000100100000100100000010000010011010001010100000111000000010000010001000000000101000000011000100100001010001001000010111010000001001000000000001010100101000101110010000100101000001000000000000011000010010001010001000000000000000100000000010000010000000000000100000110001010000101000001010110000000000100010000000100001001000000000100000011001000100000000000000100001000011000100000100000001100100000000010100000001010101001000001100010000000000100001100100000000010000000000100000100101000100000000000001000000000100010010000001001000000000000000010000010010000000000101000010101101001000101000000100000000000100000100000000000010001010000000000000010001000000000011000000000000000011000000101000000000100000000100100010001000010000000100000000000001010000000010001001100000010101010100000000000001000000010000000000000000010000101100100010001000111011000011000010000000010100100110010101000000001010000000000111100001100000000100000000000000110000000001010000010000100001000000000010101000000001001100100011000000000000000110000000011000000001000000011001100010000000010010000000011010100000000010000000000000000100000101000010001001001000000000000000000000010000000001100000000001000101000000000010010000001001000000000001101001000010011100100001000000000100001000010001001000110000000101010000000000001000110000000010001001010100001000000000100010010000111000000010000010010100000001010000110000001100000000111000000000000000000000000000100001000010010011011010100010010001101000000101000110001100010000001010001000110110001000001000110000000000010001100001010010100000100000010001000101010000000100100000000001011011000100000000010010010001010110000100100011000000010000110000000001000001110001100000001010000011010101100010000010110000000000101110000001000000000010001101000001001001001000011000001000001100000000001011101000011010000000100110000000001000110000000100000000000001010000010100001000101001110001000100001100010100000010011010000000100000001000100001000010000000000101111101100010001001100001000000000000000000101000001000011000100000000001011101101000011010001000001000000001000000110110001001010100010001000100000101000000000010000000110000011010001000000110010000000001010101000000110000110001000000100100000000100000010000000000000100000000000010000100100000100000100001000101110101010001000000000010000000010010110100011100010100000101001011000000001001100000001101001000011010001000000110000001100010001100000100000011000000000010000001110100110100000000001100010001011000100000010010010010000000101000110010000100000000010001100001010001001000000000000110010000001100000000000010000101001000000001010000010000100000001000000000001100000001100010000101000000100000001000001001010100010101110000110010000001001000001001001000001011010100000000000011011011000000100000001101001100011010000000101000000000010011000000000010000001000000000000000011000000100000001000100001110011000011001000001001001001100100000101000000000000000000000100100010010000010010100000000001001010110000100000100000000100011101011100000000000000000000000000001001000001011001001001000010000010011000010101100100110000000000000000001110011011000000110010100000010101000001100000000010000000001000000100100001000110100000000011010000000110010010000000001010001001010010000000010010111110100000000010010100000100000000100001000000111000001000000000010100000000011000010000000010000010101100000101110000001100000110010001000010000100100100000000001000011010000100001001001000000010010100101001000100011110000000110001000001100010100100000101000011101110000000001000001100000001000000000011010011000101101000001001010101101100101000010100001000010000000001010000000000101000000011010000011000110010100010000000010011010101101001000000000101001000010001100111001100001110000001000000000011000011000001000000010100101000000000010100001110010100000010000000100000100100000010000010000000111100000001000101001001000001010100110100000100000010001100000000000001010000000010001101011000001000100001110000000010110010000000101100101010000001010010101100100001001001100000100001101011000100000010000000111001000010100011010000000111101010100000000001000100011010000110001110000000110110001010000000001000110000101100000010000000001100110011001011011111111000111101100011010001000111000110100000000101001000100001001000000001010100000000001001100000101000010001000000001000000010001000000010000110000011001010100101100000001111000000000000101000100010000000010010000100000010001000010100000010000001001000111000101100111101000011001011100111100000100000010000110000100110011100011010110000100001001000001010010000010000000000101000000000001010100100010000000011011000000110100011011000000100011100000010001000010000001101000000010000000000001000010000001110011110010000000100001100000001100000010010100000110000010010000110000000010010000111111000100011110011010011011000000000000000000001100110100000100100101100001100011110001000100100001010010010001000001001011001000001010101001100100010001000000000010101110010011010110001001001100000011100000110000110011011001100000101000110000010000000010010000000001000010000011001100011101000110000011000001110010110010000000110001010001110000000111100101001101011000001000011110111001000000101010110011000000000111001100000000101001001010010000101000000110000001100100010000000000101000110000100100111010000000000101010101010100001010100010100010000000010000000001100000000000001011000000010001000100010000101101000001000011000110010000000100010000000000001011000010000001100001000010000000100100010010001110000100000001100000000010110001101010000001001010101011000000000010011010010010011010000010001011010100011000000001000100101010000000100010001011000000010110100110000110001110110001101110111000001000110010000000100000011011100010101011000110011000001010010100001001010000011000100101100101111111000110001100101001011010100100001000000001011010000100000000101110101000000010110100110000000110101100011110000100011101001010011111000101001001100001110000100001001000100010110101000010000111101110110101001000100111010010000000110111000100001000010010111001101000110001011010011110011000000010011000000000000111100000100000010000001010111110010010010010100001000100010100110001000001100000001000110100010101000000000111000111110011010110001100011011001000010001100010000011000110000100100101101110100000100000100010010001000101100110000010000011100001010011000101011111001000110001001111000100010110000000001000100011111110100101001100001100001000000111101000010000000000000110000011010001000000000100101010010000010000101000010001101111001101000010000001000110101100111000001101100101100000000011001110000101110000111000000010110001100000110010100010100000001011000011000000100001001000000000011100100001000000000100000011100000001110100100000100010010011110000101000000000100100101000100000010000010001100010100000101110010000000000001000010001101100001001000101101010010010000011011100001110000001000011001110110000100110000000110100101101101101100100001000010100001100001010100011000111010000100001010001100000000011000010000000101010001000010000010001000000001001001000010001010000010000110101000111110101001001001010001001110001010010011000001000001110000000101110000011010001001111000100100000000001100001001110000110000000010011011000100111000010001000001111110001011001000001000000000110000000000101110011000000100100100000111110000111000100000111000010110110000111110101101101101100100000010010001001101000100010011110000101010000111000000100010100100110010000000000000101110001010000000101100010110010110000010001011001010100000001010010000011110000110011010000100111010010110000000010000001011101001101000000101000101001111010001011000000011110000001000001001110011111000000110000000101100010011010001000001000000101011010011000010010000011001000001001011000010110111100100011000000001100101011001010100000110010000100100010000011111010000101111111010000010110111011110001100101101011111000011000111100001110000110001000010110000000010001000011111110110010001110100101100110010110110011001000011101110010010000000010000001010001001100011010001010001001000000110000000110011100000101001100001000001101110101110000111110011010110000001010001001000100101111000000010110101001111010000000000010011000011000000001110101111000001100000010111000011011100001100010001100000100111010000010011011010001110110110100000000100001001011110000000110011100000000100000100101101111000110000011100011101001000001011111110000100110000000001010010100010000011001100110011110100000000111000000010010100011000010100110110000101010101100000111110011101000011000110010001101000001001000100100001101000100000110110110110000100001000111001011110110000011011100000011010110101110001001000011000011000010100001010100000001111101001000001010011001100110011101010000010000100000011010001110100010000000100011101100111001011001101100100000101100100011000001000010000100110000011010001001001000000000010110110001001000100111101000000111100010010101000010001100100000000001000011010100000010010010101000011000100001011010101110010100010100110011100000101010000110110000101001100010000011011100111000000101001111000001111011110111010001000011001000110011000000000110110101100011111100011100000010101000110100000000001010000111011110001110000110010010110011011011110111000101110100100111100011100000010101010010100001001010011000001010001101100100011000000110111000011001110000100100010100011111111001111011110101110011000101101101100010010001111001001110101111111110000001111001111111110001001000001101110100010000011000110110110011100101001001010111110100101000101000100111110101011011011101101101000001000100110010001111001011001101110111010100100001011010011001000100010000100101010001010010011011101100000000000011101000111100010100001100101001000100101001010010010111101010110000001101011100101010001011011110101111010000111000100100001001111111110001000000010111000110111111101110000000110001011000000101011011001011111111111010100001111111000001000111111000111010000011010110000000010010110110011010001101010000111011001011001001100011110100110000110010001110110100101101110100010101101100010000001001110101000101101011011010001101111110000000011010111111100000100101101011110011010011010000101001010010000010101110110110000100001000110100001001111010100010011110000111010000010000001101000110001010100100100001101000011000011111011010110011010110100100100001010010000100100110010111110010100101111001110000111100101101011011110110101000010010000110100110101100000110100101010100111100010000000000001010011001000100001000000101111001010001111001001111101100001001100010010011110100010001101100100000111101010101100100100101000010010100000101011100101010110000100100100110000010010000101101001110000111001011011000110101111001111001011110100101010010000000010011101110011001101101001000110110110010110011001100110000010000000000000000010111000100110100110111110101001101001001000100111001101111010011010111011001010001010100100011001100001010010101010010010011110000000010000101100010011011110111101000000110000101101010000000001000001101101100010110000101010100000011100011000111111101000101100100001101010101001010000101100110100110011100001010000010010100010001100100000000011111011000000000011000010001011001101010111001101000000001100010101110100010111111001011100100010101000101000101010001101000110000110001000001100010010010110101100100111101100100110100111001011000101001101111000011101011010110110011101000000110000011011010101100000011100010100001010001011110001010000000001011100110100110110011001001011000011001101100000100011010001010101100011000110101101100010011010110100000110011111001010011000111011111010101100101010111100101000000100011000000001111000100101000000110101010010111000111001000001000010110101011100011100101101010101001011110000000110001010000;
		data3[16383:0] = 16384'b0000001000000000100000000100001000100101000100000000001000000010000000001000000000000000000110000000000010000000000000000000000000000000000001100000000000001000000001100001000000000000000000010000000100000000001010000000100000010000000010000000000010000000000100001000100000000000000000000010000000000010000000000000000000000000000001000000000000000001000000000000000000100000000010000000101000000000000010000000000000000000000001000001000000010010001000000000000000000000000100001000000000000000000000000100000000000000010000000000000100000001000101000000000000000010000100001000010000000000001001000000000000010000000000000000000000000000001100100001000000000000000000000000010000000000000000010000100100010000000000000000001000000000000000000000000000000000001000000000001000000100000000010101000100000000100001100100000000001000000101000001000000000000100001000100100001000001000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000001001100000000000100000000000000100000100000000000000000000011001000000000110000000000000000011100000000000000000000010000000000001000000001000000000000000000000000000000000001000000000000000000001010000000011000000000000000000000000000000000010000010000000100000000000000000000001000000001000010000000000001000001010000000000100000010000001000100000000000000000000000000000100010010000000000000000000000000010000000000001000000000000001000000000000000000001010101000010000000000000000000110000000000010000011100101000000001010000000000000010100100000000000100000000000001000010000001000000001000000000000000010000000000000010000000000000000000000000000011010000000001000000000000100000000000000000000000000000000100000000000000000100001000100000000000001000010000001010010100000100000010000100000000001001000000000000000000011000010100000001000000000000000000000000010000000000000000000100010001000000001000000000001000010000000000000000000000000000000001000000000000011000011000000000001000000000000001100000000001000000101010000000000000000000100010000010000000000010001011000010001000000000000000000000000000000110010000010100000100000000100000000000000001010000000000000001001100000000000011100011100000001000100000000000111111110001000000000100001000000100000001010000000000100000001000000000000001100000000001001100001110000001001000010000010000000000010001100000000011001000010010001000000010000000001000000000000000010010100000000000010000000000000101000000100111000100000001000000100010001100000101000000001000000001000101000000000000100000010000110000010000000100000100000000000100000100011110011000000000000010001000011001000001100000001000000000001000000000000000000000000000000001010000001000000011000000000100000000100010000000110000000000000000000000000100000000001000000000000001000000000000001001000000001000011000100000010000000000000000000000000010001000011011100100001000100001000101000000000001000000000101100000000100000000000110001000000000001000001110010001001000001000000000000000000000000000010000001000000000000100000000000000000010000010100000001000011000000000010100100000000000000100100001000001000000000000010000010000000000000000100000000000000000100000001000100000000011000110010100100000010100000000000100011000000010110000010001000000000000100000000001100000000100000010001000000000000000000000010000000000010000000000000011000000000001010000100010001000000000000001110000000100000000000000000000000000000000000000000000001000000100000000010010100000000001011000010100000000010000001010000000000100010010000001000000000010000000000000000000000000010000100000000000010000000010000000000100000010100000000010000000000011000001100000100110000000010100001010000001000010000000100000010000000100101000000000000000100111000011000000000100000100000001000000000100011010010001100011000001000000000101000000000010001000000010000001000000000110000000000000100000001011110000000000001100010000010000000000001000000000000000100000000001000000000100010000000000000010000000001100000000010100100000001100000100011000100000001000000000000000000001000000000000100000001000101000010011000111101000010000001100000100001000000010010000000000000100001000000000100010010100000000100011101100010001000010011000000001000101000001000000010000010011000010010000000010000010000000000011001101000001010010010011000000000100000010000100000001000000000010100000100010010100000010000001000000110001000000000000110001100000100011000000100100000000000000000000100000001010000000000001000001010000100000011000000010010011000010000100100101001000000000100000000100100000000000000000000100100000000000001100110110000010000000001100100000101001100010000010000000100001100000000010010001000000100001000001000000011010010000010100010101000011000001000000011000000000010000001100001001000001001000100010000000000000000000000010000110000000000000000010000010000010010110110000001000100000010000000010000100001001101000000000000100000000000000000001000000000000001000000000101000000000010000001000010010100001100000000000000000000000110000100000100001000000000000000001100000000001000000100001010010000000011000000000010000110001100000011001100000000000100100100000000001011000000000100010000011000010000000100000000001000000011000010100010010000000000000000100000000000011100000000000001000110100000010000101010000000000001100100001000001000100000000000010000010100101100010000001000100100000000000100000010011010000010000000001001000000011010000011000001100000001000000000000010000011000001100000000000000000100000001110000100010001000000010101011000001000000100100100110001000000000000000100001110110000000010010101001011001101000000000010000000000100100100100001000001000010000010000001000001000000010000000000101010110100010001010000001010010000011000000101101000000000010011000000010000000000100000101000100000010010000101000000000000001000001000001000000100001000000000110010000000001100100000000010100000010001010000011100000000100100001000000000000000010000001000100000110000001000100000000010100000000001100000001000000100000000010000000000000000000000000000010001000010010000000001000100101000001000000000001000010001001110001001011000001011010101110001011001000100000000000000100001000000101000000000010000100000000101000000000100010000100010000000101100100000100101100111000000000000010001001010000000101010000010000001111001010111110001000001001000001000001000010110000101010011000001001000010001000110000100010100000000000000000101100000000000000100111000110001101101100110000000000000000000100001000001000000000000001010000000000100000000100000001010000100000011100001000010110000000000100010100001011100000100010000001010110001010001001000001000101000100100001111000000000101010000100000010100001000011101010011000000000100000000011000000010001000100100000000011000110000001000100010000000101010100000001000100000000000001010100000000010010000010010010001000000010011000000111001100101100000001110000110001000000000001100100000100100000100010010000010000001000100010000000000000110010100110000100000111000100000000010001000000000000011000010000100001000000000000101001100010010101000000010000100110010001000100100000000000001001001000000000101001100001100000000100000010001000000000111001001000000000000001000100000000000110011111010010000000000000000001100000010000000000000001000000000001100001100000101000010111100000100000011011010000000000000000000010000010001110001011000000000000000100001001000011000000100010000001110110000000000000001000100001000001000101001000000110011011001000000001000000010000100001010001000110101000100000010000000000000110000000000111000000010101000000000000000000010010001010010011011000100100100001111001000000000001010000000000111010010000000000100000010001000000000000010000000001000000000000001000000101001010001000000011110000110101000001100100001000000000011010000110000000000100000111000001000001110111000000000000010000001001001000000000000011010100100000010001001110100000100001000001000000000000000000100110000100000001000000001000000100011000001000000010100000010111000001010001000000001000101000010000010101000000000000001000000000000001100110101001011100000000000111000010101010000000011010001000000010001000010000001111101001000010000101011000000001010011001000101000100001000101001001000100001001110000010100001001000010000100100000001100111010001011100101010001000010101010000001001010000011010000001001000011011100011000100010001000100100000100000000010100010110000001000001010001011010000110100001001000011101000001100011100101001010101110001100011011011010010001001100100100000100001000101000001100000000000000000010001000010000001100110010001000011001000110000010111000110110001100101000000000000100100001010010010010000000110001000001100100100110100111010000110000001100000010001100000110001010001000001000100000100001110011001100001010101000100000110000011010001110000000000000000100011000110010000101001100010001101001010010010000001100010010101010000000100001011100000100010010101100010100100001100000011001101000000100000101000001001000100000010000010011000001001110001010011000010100010000011101000010000011101111100001101010001011100001100010000010000100110001011011000000001010100010001101000110001000011001001000000000100101011000111100000000100100010000001100000000000010001100001101001000010001001000110010000001100011000000111001001100000000010000100101001000001110000010001101000001011001010000001000000001100001010011001110000001100000000000100010000100000100000010010100100000001000000000010011011000001001011000011111100000110110001000010000011101000000111101100100001000111110001000010000010100000011010000100001000001010001001000100000010010100010100000000100000100110101010010000000000001000000101011010000101000101110100010001100000000000010101010001000000101001000000000100001110100000001101100110000010101010100010011001101101011001100000000100001001110100000010000110000101001000001000100000000000000101100000101010110010010000011000000000000000000100000000001011000000000101000001001110000100010000000110001001000011110001100000100110101111010000000010100100101000100100010001011001110001000100000000111011001000000000100100011000101000101111000100010100000010000110011001001100000000011100001000000011000000100000000100100000010100000100011110000100000111101010110000000000100101000100001100010001010100001001011000010101000100010110001111101000111010000101000010011110100000001010101001101101000010001010000101110010000000100000100011110100001100100010000000001000001100000000010010001101110101101100011000101011001000100000100000001000000010000000010000001001000001101001010011010010001001000011000100000000010000000010000000110101001001010001000001000001000000110101000000000110011100100001001000000000001000101100001000100001100000000000000100001111010000100011111001100000000110010100111100101001100101111001000100011000001000110001010001100011001001101000000001010100000000010101101000000100010001100010010011100010000010101011111101001101001110010000110111000100100111001111011000001001100010100100101000011110000001000100100110110000010000000010010000010010100010010001010110100010000011100111000110011000001101111111001010000101000000001111111010001101011101010000000101001011100001111001100011000000010100000110101100101111001110111001110100100010101110110001100000100100010000010000110010101100001111011001100000000110011101100000110000110001001100011000110100101100001000000010110011010000000000000100100101000000101011001010011110000001011000110110010001100010010000100011001010010010100001010110111100010000000100011011011000001110111010000010101011001001110101010101000001101001101100000000010001100001110010010011110101010010010010111000100010000000000001000001100110110000010010000001110100110001001010001000010000000100000101001110100001001000001010001111100000110000100000000001100110000001010100110000001000000101100100011010100000000100000110110001001000110110111111111100000110100000101011101000100000111100110000100000111000001100111101000001110101000010111001100110000000111000000001010000100010011001000010001100001001110010001000100000000100001010100010010010110110000001101010000000111100001101111001101010010001001100000001000010001111001001100000001000110110001100100010011000000111001011000011000000011000000111000101100011000001000001100001000110110001101110010001000000000011110010101011101000001000101011011000100001000100000000101001001111111010000011010100000101000101010000010011101100010111000100010000001001010100100100111100100011111000000011001101100110001111100010100111000010010010111011001101101010000011000001000010000000001110100011100110111000001001010101110001000000110000101000001000011110111010010000011100010000001101001001100011011100000000101100001000110101010100000111010100011000111001000001110100111001000000010010101100000001100000000011110101001111001111011001000000001001010001010000101011001010100001100000001000001010011000001000010101011001101100100001010010100001010011001011000001011101100111010010011010010100010001011101011000010100100000000101001001011100110100101001010110100010101101101100100000100101101100111001111011000010100001001110110100001011111011000000000111110101010111011000000010000011101000110000001000000110011000100010011010010011101000000110000010001011001010000100010010011000010110000001011000101100001010001010010011001100110101011110011100100001000000000101110010000000101100101001100110010110010001100001100000110110000000100011001000000100000000111101100000000000010100101111110110010101110010000101000100001101001000000001001101010101001001001001000000111110000110011010111010110100000001110000000000000110001100010110011010100001010011101000011000010010111000010001101001010000000100000001011101000000000001001001101110110001101100000110000100001011001011000010111000011011000110110100001100010010000100010111001110010010001101001000111011000110101011101000100001100110101100001100001100011101011000010010110000000011010110101101010111001100101101001000000111000000010010100001100010001000111111100101000011010001011010000000010000000011010010111100000110010110101000000001110111000000111001100111010011011101011011110100011011010100000011001010001110000111001100010100010000010100001110001100001010000110010001011001001100000001011110110001111010101000000011000011000110000111010000000010000000111000011110100000000000011000000000011010100110010110000000100010001111000000000100100110100010000111010001001000001110010000001101010000101000010000000111100111110001001010111100100101000101010010111010100011010111101101010001010001011010001011000001110001001101010000010011001100001111101000010101010001010101100000011000010001110000001000100011101011001001001110000111110011000001100100110010101000001001101000010100100000000110101110001010100001101000000110101010100111110000101110000000110001010011101101010100000000010000011001101111100101101000010010011110000010000010110111111110011111001011001011011110001000010000001011110001101100110110011111100100000101100001110111011101011001010110000010000101001100110101011011001011010100110001011111001100001111001110000001100000011100010000000010000111001001000001001100100001011011001101001101000110101010010111100110100000101000010011011110101010001011101000011010000110010010110000000000010000000101101100011100000000011001110100111010000100101011111111001000111001000001110011011110011000011101110110010000100011110011101100100010011001010101111011010101100100001010010001110111010001011110110100110101100010111100010111000010000100111100010110001101000001001100111101100100010011010101001100101111000001011111000001001000010010011001000111101010011010001001010100000000010010001110110100001010001010110100111001110101010101010010000010111010101111000100110001110010110001000110011101100011011111000111000101011011101001000100111010001001000011111110010111111100010100100100100010100001111101100111011000101100100000011000110011111100111000101010101010100010100010010110001101000100011110110000101010001000110011101100010100110110111111011000000000000011000100111101010110010011001000110101010101010101001010000101001110010001001000011000100100100100101001100100000011100000000001000000110001010101011011001101110010000110001001010000100111110011100100000110101011011001000000000001010100011001000101010011110010111111010000010110010100110001101001110001100011001100000000011000100011111010100000010100010000000100011011011100;
		started = 1'b0;
		num[14:0] <= 15'b0;
		startlast <= 1'b1;
		show0[6:0] <= 7'b1111111; // 左边
		show1[6:0] <= 7'b1111111;
		show2[6:0] <= 7'b1111111;
		show3[6:0] <= 7'b1111111;
		show4[6:0] <= 7'b1111111;
		show5[6:0] <= 7'b1111111;
		score[11:0] <= 12'b0;
		LED[7:0] <= 8'b0;
		failed <= 0;
	end

	always@(posedge clk)
	begin
		// start
		if(!start && startlast)
		begin
			score = 0;
			num <= 32 * {switch[5:0]};
			started <= 1;
				show0[6:0] <= 7'b1111111; // 左边
		show1[6:0] <= 7'b1111111;
		show2[6:0] <= 7'b1111111;
		show3[6:0] <= 7'b1111111;
		show4[6:0] <= 7'b1111111;
		show5[6:0] <= 7'b1111111;
			button0Last = 1;
			button1Last = 1;
			button2Last = 1;
		end
		startlast <= start;

		// cleared the item
		if(!button[2:2] && button2Last)
			begin
				if(show0[3:3]==0)
				begin
					score = score + 1;
					show0[3:3] <= 1;
				end
				else
				begin
					if(show1[3:3]==0)
					begin
						score = score + 1;
						show1[3:3] <= 1;
					end
					else
						failed <= 1;
				end
			end
		if(!button[0:0] && button0Last)
			begin
				if(show0[6:6]==0)
				begin
					score = score + 1;
					show0[6:6] <= 1;
				end
				else
				begin
					if(show1[6:6]==0)
					begin
						score = score + 1;
						show1[6:6] <= 1;
					end
					else
						failed <= 1;
				end
			end
		if(!button[1:1] && button1Last)
			begin
			if(show0[0:0]==0)
				begin
					score = score + 1;
					show0[0:0] <= 1;
				end
				else
				begin
					if(show1[0:0]==0)
					begin
						score = score + 1;
						show1[0:0] <= 1;
					end
					else
						failed <= 1;
				end
			end
			button0Last = button[0:0];
			button1Last = button[1:1];
			button2Last = button[2:2];
		// record now times
		state[10:0] <= state[10:0] + 1;
		if(started)
		begin
			// if time counted 500 * speed (ms)
			if(state[10:0] > (speed[1:0] + 2'b01) * 500)
			begin
					 LED = LED + 1;
				num <= num + 1;
				if(num > 2047)
					num <= 0;
				state[10:0] <= 11'b0;
				if(show0[6:6] == 0 || show0[3:3] == 0 || show0[0:0] == 0 || failed)
				begin
							failed <= 0;
					LED = 0;
					started <= 0;
					// 显示得分，得分清零
					// show0-5
					//读出个位
					out = score % 10;
					case (out)
						4'b0000:{show5}<=7'b0000001;	//0
						4'b0001:{show5}<=7'b1001111;	//1
						4'b0010:{show5}<=7'b0010010;	//2
						4'b0011:{show5}<=7'b0000110;	//3
						4'b0100:{show5}<=7'b1001100;	//4
						4'b0101:{show5}<=7'b0100100;	//5
						4'b0110:{show5}<=7'b0100000;	//6
						4'b0111:{show5}<=7'b0001111;	//7
						4'b1000:{show5}<=7'b0000000;	//8
						4'b1001:{show5}<=7'b0000100;	//9
					endcase
					score = score / 10;
					out = score % 10;
					//读出十位
					case (out)
						4'b0000:{show4}<=7'b0000001;	//0
						4'b0001:{show4}<=7'b1001111;	//1
						4'b0010:{show4}<=7'b0010010;	//2
						4'b0011:{show4}<=7'b0000110;	//3
						4'b0100:{show4}<=7'b1001100;	//4
						4'b0101:{show4}<=7'b0100100;	//5
						4'b0110:{show4}<=7'b0100000;	//6
						4'b0111:{show4}<=7'b0001111;	//7
						4'b1000:{show4}<=7'b0000000;	//8
						4'b1001:{show4}<=7'b0000100;	//9
					endcase
					score = score / 10;
					out = score % 10;
					//读出百位
					case (out)
						4'b0000:{show3}<=7'b0000001;	//0
						4'b0001:{show3}<=7'b1001111;	//1
						4'b0010:{show3}<=7'b0010010;	//2
						4'b0011:{show3}<=7'b0000110;	//3
						4'b0100:{show3}<=7'b1001100;	//4
						4'b0101:{show3}<=7'b0100100;	//5
						4'b0110:{show3}<=7'b0100000;	//6
						4'b0111:{show3}<=7'b0001111;	//7
						4'b1000:{show3}<=7'b0000000;	//8
						4'b1001:{show3}<=7'b0000100;	//9
					endcase
					score = score / 10;
					out = score % 10;
					//读出千位
					case (out)
						4'b0000:{show2}<=7'b0000001;	//0
						4'b0001:{show2}<=7'b1001111;	//1
						4'b0010:{show2}<=7'b0010010;	//2
						4'b0011:{show2}<=7'b0000110;	//3
						4'b0100:{show2}<=7'b1001100;	//4
						4'b0101:{show2}<=7'b0100100;	//5
						4'b0110:{show2}<=7'b0100000;	//6
						4'b0111:{show2}<=7'b0001111;	//7
						4'b1000:{show2}<=7'b0000000;	//8
						4'b1001:{show2}<=7'b0000100;	//9
					endcase
					{show1}<=7'b1111111;
					{show0}<=7'b1001000;
					score = 0;
				end
					else
					begin
                case(num)
                    0:
                        begin
                        left <= data1[0:0];
                            middle <= data2[0:0];
                            right <= data3[0:0];
                        end
                    1:
                        begin
                        left <= data1[1:1];
                            middle <= data2[1:1];
                            right <= data3[1:1];
                        end
                    2:
                        begin
                        left <= data1[2:2];
                            middle <= data2[2:2];
                            right <= data3[2:2];
                        end
                    3:
                        begin
                        left <= data1[3:3];
                            middle <= data2[3:3];
                            right <= data3[3:3];
                        end
                    4:
                        begin
                        left <= data1[4:4];
                            middle <= data2[4:4];
                            right <= data3[4:4];
                        end
                    5:
                        begin
                        left <= data1[5:5];
                            middle <= data2[5:5];
                            right <= data3[5:5];
                        end
                    6:
                        begin
                        left <= data1[6:6];
                            middle <= data2[6:6];
                            right <= data3[6:6];
                        end
                    7:
                        begin
                        left <= data1[7:7];
                            middle <= data2[7:7];
                            right <= data3[7:7];
                        end
                    8:
                        begin
                        left <= data1[8:8];
                            middle <= data2[8:8];
                            right <= data3[8:8];
                        end
                    9:
                        begin
                        left <= data1[9:9];
                            middle <= data2[9:9];
                            right <= data3[9:9];
                        end
                    10:
                        begin
                        left <= data1[10:10];
                            middle <= data2[10:10];
                            right <= data3[10:10];
                        end
                    11:
                        begin
                        left <= data1[11:11];
                            middle <= data2[11:11];
                            right <= data3[11:11];
                        end
                    12:
                        begin
                        left <= data1[12:12];
                            middle <= data2[12:12];
                            right <= data3[12:12];
                        end
                    13:
                        begin
                        left <= data1[13:13];
                            middle <= data2[13:13];
                            right <= data3[13:13];
                        end
                    14:
                        begin
                        left <= data1[14:14];
                            middle <= data2[14:14];
                            right <= data3[14:14];
                        end
                    15:
                        begin
                        left <= data1[15:15];
                            middle <= data2[15:15];
                            right <= data3[15:15];
                        end
                    16:
                        begin
                        left <= data1[16:16];
                            middle <= data2[16:16];
                            right <= data3[16:16];
                        end
                    17:
                        begin
                        left <= data1[17:17];
                            middle <= data2[17:17];
                            right <= data3[17:17];
                        end
                    18:
                        begin
                        left <= data1[18:18];
                            middle <= data2[18:18];
                            right <= data3[18:18];
                        end
                    19:
                        begin
                        left <= data1[19:19];
                            middle <= data2[19:19];
                            right <= data3[19:19];
                        end
                    20:
                        begin
                        left <= data1[20:20];
                            middle <= data2[20:20];
                            right <= data3[20:20];
                        end
                    21:
                        begin
                        left <= data1[21:21];
                            middle <= data2[21:21];
                            right <= data3[21:21];
                        end
                    22:
                        begin
                        left <= data1[22:22];
                            middle <= data2[22:22];
                            right <= data3[22:22];
                        end
                    23:
                        begin
                        left <= data1[23:23];
                            middle <= data2[23:23];
                            right <= data3[23:23];
                        end
                    24:
                        begin
                        left <= data1[24:24];
                            middle <= data2[24:24];
                            right <= data3[24:24];
                        end
                    25:
                        begin
                        left <= data1[25:25];
                            middle <= data2[25:25];
                            right <= data3[25:25];
                        end
                    26:
                        begin
                        left <= data1[26:26];
                            middle <= data2[26:26];
                            right <= data3[26:26];
                        end
                    27:
                        begin
                        left <= data1[27:27];
                            middle <= data2[27:27];
                            right <= data3[27:27];
                        end
                    28:
                        begin
                        left <= data1[28:28];
                            middle <= data2[28:28];
                            right <= data3[28:28];
                        end
                    29:
                        begin
                        left <= data1[29:29];
                            middle <= data2[29:29];
                            right <= data3[29:29];
                        end
                    30:
                        begin
                        left <= data1[30:30];
                            middle <= data2[30:30];
                            right <= data3[30:30];
                        end
                    31:
                        begin
                        left <= data1[31:31];
                            middle <= data2[31:31];
                            right <= data3[31:31];
                        end
                    32:
                        begin
                        left <= data1[32:32];
                            middle <= data2[32:32];
                            right <= data3[32:32];
                        end
                    33:
                        begin
                        left <= data1[33:33];
                            middle <= data2[33:33];
                            right <= data3[33:33];
                        end
                    34:
                        begin
                        left <= data1[34:34];
                            middle <= data2[34:34];
                            right <= data3[34:34];
                        end
                    35:
                        begin
                        left <= data1[35:35];
                            middle <= data2[35:35];
                            right <= data3[35:35];
                        end
                    36:
                        begin
                        left <= data1[36:36];
                            middle <= data2[36:36];
                            right <= data3[36:36];
                        end
                    37:
                        begin
                        left <= data1[37:37];
                            middle <= data2[37:37];
                            right <= data3[37:37];
                        end
                    38:
                        begin
                        left <= data1[38:38];
                            middle <= data2[38:38];
                            right <= data3[38:38];
                        end
                    39:
                        begin
                        left <= data1[39:39];
                            middle <= data2[39:39];
                            right <= data3[39:39];
                        end
                    40:
                        begin
                        left <= data1[40:40];
                            middle <= data2[40:40];
                            right <= data3[40:40];
                        end
                    41:
                        begin
                        left <= data1[41:41];
                            middle <= data2[41:41];
                            right <= data3[41:41];
                        end
                    42:
                        begin
                        left <= data1[42:42];
                            middle <= data2[42:42];
                            right <= data3[42:42];
                        end
                    43:
                        begin
                        left <= data1[43:43];
                            middle <= data2[43:43];
                            right <= data3[43:43];
                        end
                    44:
                        begin
                        left <= data1[44:44];
                            middle <= data2[44:44];
                            right <= data3[44:44];
                        end
                    45:
                        begin
                        left <= data1[45:45];
                            middle <= data2[45:45];
                            right <= data3[45:45];
                        end
                    46:
                        begin
                        left <= data1[46:46];
                            middle <= data2[46:46];
                            right <= data3[46:46];
                        end
                    47:
                        begin
                        left <= data1[47:47];
                            middle <= data2[47:47];
                            right <= data3[47:47];
                        end
                    48:
                        begin
                        left <= data1[48:48];
                            middle <= data2[48:48];
                            right <= data3[48:48];
                        end
                    49:
                        begin
                        left <= data1[49:49];
                            middle <= data2[49:49];
                            right <= data3[49:49];
                        end
                    50:
                        begin
                        left <= data1[50:50];
                            middle <= data2[50:50];
                            right <= data3[50:50];
                        end
                    51:
                        begin
                        left <= data1[51:51];
                            middle <= data2[51:51];
                            right <= data3[51:51];
                        end
                    52:
                        begin
                        left <= data1[52:52];
                            middle <= data2[52:52];
                            right <= data3[52:52];
                        end
                    53:
                        begin
                        left <= data1[53:53];
                            middle <= data2[53:53];
                            right <= data3[53:53];
                        end
                    54:
                        begin
                        left <= data1[54:54];
                            middle <= data2[54:54];
                            right <= data3[54:54];
                        end
                    55:
                        begin
                        left <= data1[55:55];
                            middle <= data2[55:55];
                            right <= data3[55:55];
                        end
                    56:
                        begin
                        left <= data1[56:56];
                            middle <= data2[56:56];
                            right <= data3[56:56];
                        end
                    57:
                        begin
                        left <= data1[57:57];
                            middle <= data2[57:57];
                            right <= data3[57:57];
                        end
                    58:
                        begin
                        left <= data1[58:58];
                            middle <= data2[58:58];
                            right <= data3[58:58];
                        end
                    59:
                        begin
                        left <= data1[59:59];
                            middle <= data2[59:59];
                            right <= data3[59:59];
                        end
                    60:
                        begin
                        left <= data1[60:60];
                            middle <= data2[60:60];
                            right <= data3[60:60];
                        end
                    61:
                        begin
                        left <= data1[61:61];
                            middle <= data2[61:61];
                            right <= data3[61:61];
                        end
                    62:
                        begin
                        left <= data1[62:62];
                            middle <= data2[62:62];
                            right <= data3[62:62];
                        end
                    63:
                        begin
                        left <= data1[63:63];
                            middle <= data2[63:63];
                            right <= data3[63:63];
                        end
                    64:
                        begin
                        left <= data1[64:64];
                            middle <= data2[64:64];
                            right <= data3[64:64];
                        end
                    65:
                        begin
                        left <= data1[65:65];
                            middle <= data2[65:65];
                            right <= data3[65:65];
                        end
                    66:
                        begin
                        left <= data1[66:66];
                            middle <= data2[66:66];
                            right <= data3[66:66];
                        end
                    67:
                        begin
                        left <= data1[67:67];
                            middle <= data2[67:67];
                            right <= data3[67:67];
                        end
                    68:
                        begin
                        left <= data1[68:68];
                            middle <= data2[68:68];
                            right <= data3[68:68];
                        end
                    69:
                        begin
                        left <= data1[69:69];
                            middle <= data2[69:69];
                            right <= data3[69:69];
                        end
                    70:
                        begin
                        left <= data1[70:70];
                            middle <= data2[70:70];
                            right <= data3[70:70];
                        end
                    71:
                        begin
                        left <= data1[71:71];
                            middle <= data2[71:71];
                            right <= data3[71:71];
                        end
                    72:
                        begin
                        left <= data1[72:72];
                            middle <= data2[72:72];
                            right <= data3[72:72];
                        end
                    73:
                        begin
                        left <= data1[73:73];
                            middle <= data2[73:73];
                            right <= data3[73:73];
                        end
                    74:
                        begin
                        left <= data1[74:74];
                            middle <= data2[74:74];
                            right <= data3[74:74];
                        end
                    75:
                        begin
                        left <= data1[75:75];
                            middle <= data2[75:75];
                            right <= data3[75:75];
                        end
                    76:
                        begin
                        left <= data1[76:76];
                            middle <= data2[76:76];
                            right <= data3[76:76];
                        end
                    77:
                        begin
                        left <= data1[77:77];
                            middle <= data2[77:77];
                            right <= data3[77:77];
                        end
                    78:
                        begin
                        left <= data1[78:78];
                            middle <= data2[78:78];
                            right <= data3[78:78];
                        end
                    79:
                        begin
                        left <= data1[79:79];
                            middle <= data2[79:79];
                            right <= data3[79:79];
                        end
                    80:
                        begin
                        left <= data1[80:80];
                            middle <= data2[80:80];
                            right <= data3[80:80];
                        end
                    81:
                        begin
                        left <= data1[81:81];
                            middle <= data2[81:81];
                            right <= data3[81:81];
                        end
                    82:
                        begin
                        left <= data1[82:82];
                            middle <= data2[82:82];
                            right <= data3[82:82];
                        end
                    83:
                        begin
                        left <= data1[83:83];
                            middle <= data2[83:83];
                            right <= data3[83:83];
                        end
                    84:
                        begin
                        left <= data1[84:84];
                            middle <= data2[84:84];
                            right <= data3[84:84];
                        end
                    85:
                        begin
                        left <= data1[85:85];
                            middle <= data2[85:85];
                            right <= data3[85:85];
                        end
                    86:
                        begin
                        left <= data1[86:86];
                            middle <= data2[86:86];
                            right <= data3[86:86];
                        end
                    87:
                        begin
                        left <= data1[87:87];
                            middle <= data2[87:87];
                            right <= data3[87:87];
                        end
                    88:
                        begin
                        left <= data1[88:88];
                            middle <= data2[88:88];
                            right <= data3[88:88];
                        end
                    89:
                        begin
                        left <= data1[89:89];
                            middle <= data2[89:89];
                            right <= data3[89:89];
                        end
                    90:
                        begin
                        left <= data1[90:90];
                            middle <= data2[90:90];
                            right <= data3[90:90];
                        end
                    91:
                        begin
                        left <= data1[91:91];
                            middle <= data2[91:91];
                            right <= data3[91:91];
                        end
                    92:
                        begin
                        left <= data1[92:92];
                            middle <= data2[92:92];
                            right <= data3[92:92];
                        end
                    93:
                        begin
                        left <= data1[93:93];
                            middle <= data2[93:93];
                            right <= data3[93:93];
                        end
                    94:
                        begin
                        left <= data1[94:94];
                            middle <= data2[94:94];
                            right <= data3[94:94];
                        end
                    95:
                        begin
                        left <= data1[95:95];
                            middle <= data2[95:95];
                            right <= data3[95:95];
                        end
                    96:
                        begin
                        left <= data1[96:96];
                            middle <= data2[96:96];
                            right <= data3[96:96];
                        end
                    97:
                        begin
                        left <= data1[97:97];
                            middle <= data2[97:97];
                            right <= data3[97:97];
                        end
                    98:
                        begin
                        left <= data1[98:98];
                            middle <= data2[98:98];
                            right <= data3[98:98];
                        end
                    99:
                        begin
                        left <= data1[99:99];
                            middle <= data2[99:99];
                            right <= data3[99:99];
                        end
                    100:
                        begin
                        left <= data1[100:100];
                            middle <= data2[100:100];
                            right <= data3[100:100];
                        end
                    101:
                        begin
                        left <= data1[101:101];
                            middle <= data2[101:101];
                            right <= data3[101:101];
                        end
                    102:
                        begin
                        left <= data1[102:102];
                            middle <= data2[102:102];
                            right <= data3[102:102];
                        end
                    103:
                        begin
                        left <= data1[103:103];
                            middle <= data2[103:103];
                            right <= data3[103:103];
                        end
                    104:
                        begin
                        left <= data1[104:104];
                            middle <= data2[104:104];
                            right <= data3[104:104];
                        end
                    105:
                        begin
                        left <= data1[105:105];
                            middle <= data2[105:105];
                            right <= data3[105:105];
                        end
                    106:
                        begin
                        left <= data1[106:106];
                            middle <= data2[106:106];
                            right <= data3[106:106];
                        end
                    107:
                        begin
                        left <= data1[107:107];
                            middle <= data2[107:107];
                            right <= data3[107:107];
                        end
                    108:
                        begin
                        left <= data1[108:108];
                            middle <= data2[108:108];
                            right <= data3[108:108];
                        end
                    109:
                        begin
                        left <= data1[109:109];
                            middle <= data2[109:109];
                            right <= data3[109:109];
                        end
                    110:
                        begin
                        left <= data1[110:110];
                            middle <= data2[110:110];
                            right <= data3[110:110];
                        end
                    111:
                        begin
                        left <= data1[111:111];
                            middle <= data2[111:111];
                            right <= data3[111:111];
                        end
                    112:
                        begin
                        left <= data1[112:112];
                            middle <= data2[112:112];
                            right <= data3[112:112];
                        end
                    113:
                        begin
                        left <= data1[113:113];
                            middle <= data2[113:113];
                            right <= data3[113:113];
                        end
                    114:
                        begin
                        left <= data1[114:114];
                            middle <= data2[114:114];
                            right <= data3[114:114];
                        end
                    115:
                        begin
                        left <= data1[115:115];
                            middle <= data2[115:115];
                            right <= data3[115:115];
                        end
                    116:
                        begin
                        left <= data1[116:116];
                            middle <= data2[116:116];
                            right <= data3[116:116];
                        end
                    117:
                        begin
                        left <= data1[117:117];
                            middle <= data2[117:117];
                            right <= data3[117:117];
                        end
                    118:
                        begin
                        left <= data1[118:118];
                            middle <= data2[118:118];
                            right <= data3[118:118];
                        end
                    119:
                        begin
                        left <= data1[119:119];
                            middle <= data2[119:119];
                            right <= data3[119:119];
                        end
                    120:
                        begin
                        left <= data1[120:120];
                            middle <= data2[120:120];
                            right <= data3[120:120];
                        end
                    121:
                        begin
                        left <= data1[121:121];
                            middle <= data2[121:121];
                            right <= data3[121:121];
                        end
                    122:
                        begin
                        left <= data1[122:122];
                            middle <= data2[122:122];
                            right <= data3[122:122];
                        end
                    123:
                        begin
                        left <= data1[123:123];
                            middle <= data2[123:123];
                            right <= data3[123:123];
                        end
                    124:
                        begin
                        left <= data1[124:124];
                            middle <= data2[124:124];
                            right <= data3[124:124];
                        end
                    125:
                        begin
                        left <= data1[125:125];
                            middle <= data2[125:125];
                            right <= data3[125:125];
                        end
                    126:
                        begin
                        left <= data1[126:126];
                            middle <= data2[126:126];
                            right <= data3[126:126];
                        end
                    127:
                        begin
                        left <= data1[127:127];
                            middle <= data2[127:127];
                            right <= data3[127:127];
                        end
                    128:
                        begin
                        left <= data1[128:128];
                            middle <= data2[128:128];
                            right <= data3[128:128];
                        end
                    129:
                        begin
                        left <= data1[129:129];
                            middle <= data2[129:129];
                            right <= data3[129:129];
                        end
                    130:
                        begin
                        left <= data1[130:130];
                            middle <= data2[130:130];
                            right <= data3[130:130];
                        end
                    131:
                        begin
                        left <= data1[131:131];
                            middle <= data2[131:131];
                            right <= data3[131:131];
                        end
                    132:
                        begin
                        left <= data1[132:132];
                            middle <= data2[132:132];
                            right <= data3[132:132];
                        end
                    133:
                        begin
                        left <= data1[133:133];
                            middle <= data2[133:133];
                            right <= data3[133:133];
                        end
                    134:
                        begin
                        left <= data1[134:134];
                            middle <= data2[134:134];
                            right <= data3[134:134];
                        end
                    135:
                        begin
                        left <= data1[135:135];
                            middle <= data2[135:135];
                            right <= data3[135:135];
                        end
                    136:
                        begin
                        left <= data1[136:136];
                            middle <= data2[136:136];
                            right <= data3[136:136];
                        end
                    137:
                        begin
                        left <= data1[137:137];
                            middle <= data2[137:137];
                            right <= data3[137:137];
                        end
                    138:
                        begin
                        left <= data1[138:138];
                            middle <= data2[138:138];
                            right <= data3[138:138];
                        end
                    139:
                        begin
                        left <= data1[139:139];
                            middle <= data2[139:139];
                            right <= data3[139:139];
                        end
                    140:
                        begin
                        left <= data1[140:140];
                            middle <= data2[140:140];
                            right <= data3[140:140];
                        end
                    141:
                        begin
                        left <= data1[141:141];
                            middle <= data2[141:141];
                            right <= data3[141:141];
                        end
                    142:
                        begin
                        left <= data1[142:142];
                            middle <= data2[142:142];
                            right <= data3[142:142];
                        end
                    143:
                        begin
                        left <= data1[143:143];
                            middle <= data2[143:143];
                            right <= data3[143:143];
                        end
                    144:
                        begin
                        left <= data1[144:144];
                            middle <= data2[144:144];
                            right <= data3[144:144];
                        end
                    145:
                        begin
                        left <= data1[145:145];
                            middle <= data2[145:145];
                            right <= data3[145:145];
                        end
                    146:
                        begin
                        left <= data1[146:146];
                            middle <= data2[146:146];
                            right <= data3[146:146];
                        end
                    147:
                        begin
                        left <= data1[147:147];
                            middle <= data2[147:147];
                            right <= data3[147:147];
                        end
                    148:
                        begin
                        left <= data1[148:148];
                            middle <= data2[148:148];
                            right <= data3[148:148];
                        end
                    149:
                        begin
                        left <= data1[149:149];
                            middle <= data2[149:149];
                            right <= data3[149:149];
                        end
                    150:
                        begin
                        left <= data1[150:150];
                            middle <= data2[150:150];
                            right <= data3[150:150];
                        end
                    151:
                        begin
                        left <= data1[151:151];
                            middle <= data2[151:151];
                            right <= data3[151:151];
                        end
                    152:
                        begin
                        left <= data1[152:152];
                            middle <= data2[152:152];
                            right <= data3[152:152];
                        end
                    153:
                        begin
                        left <= data1[153:153];
                            middle <= data2[153:153];
                            right <= data3[153:153];
                        end
                    154:
                        begin
                        left <= data1[154:154];
                            middle <= data2[154:154];
                            right <= data3[154:154];
                        end
                    155:
                        begin
                        left <= data1[155:155];
                            middle <= data2[155:155];
                            right <= data3[155:155];
                        end
                    156:
                        begin
                        left <= data1[156:156];
                            middle <= data2[156:156];
                            right <= data3[156:156];
                        end
                    157:
                        begin
                        left <= data1[157:157];
                            middle <= data2[157:157];
                            right <= data3[157:157];
                        end
                    158:
                        begin
                        left <= data1[158:158];
                            middle <= data2[158:158];
                            right <= data3[158:158];
                        end
                    159:
                        begin
                        left <= data1[159:159];
                            middle <= data2[159:159];
                            right <= data3[159:159];
                        end
                    160:
                        begin
                        left <= data1[160:160];
                            middle <= data2[160:160];
                            right <= data3[160:160];
                        end
                    161:
                        begin
                        left <= data1[161:161];
                            middle <= data2[161:161];
                            right <= data3[161:161];
                        end
                    162:
                        begin
                        left <= data1[162:162];
                            middle <= data2[162:162];
                            right <= data3[162:162];
                        end
                    163:
                        begin
                        left <= data1[163:163];
                            middle <= data2[163:163];
                            right <= data3[163:163];
                        end
                    164:
                        begin
                        left <= data1[164:164];
                            middle <= data2[164:164];
                            right <= data3[164:164];
                        end
                    165:
                        begin
                        left <= data1[165:165];
                            middle <= data2[165:165];
                            right <= data3[165:165];
                        end
                    166:
                        begin
                        left <= data1[166:166];
                            middle <= data2[166:166];
                            right <= data3[166:166];
                        end
                    167:
                        begin
                        left <= data1[167:167];
                            middle <= data2[167:167];
                            right <= data3[167:167];
                        end
                    168:
                        begin
                        left <= data1[168:168];
                            middle <= data2[168:168];
                            right <= data3[168:168];
                        end
                    169:
                        begin
                        left <= data1[169:169];
                            middle <= data2[169:169];
                            right <= data3[169:169];
                        end
                    170:
                        begin
                        left <= data1[170:170];
                            middle <= data2[170:170];
                            right <= data3[170:170];
                        end
                    171:
                        begin
                        left <= data1[171:171];
                            middle <= data2[171:171];
                            right <= data3[171:171];
                        end
                    172:
                        begin
                        left <= data1[172:172];
                            middle <= data2[172:172];
                            right <= data3[172:172];
                        end
                    173:
                        begin
                        left <= data1[173:173];
                            middle <= data2[173:173];
                            right <= data3[173:173];
                        end
                    174:
                        begin
                        left <= data1[174:174];
                            middle <= data2[174:174];
                            right <= data3[174:174];
                        end
                    175:
                        begin
                        left <= data1[175:175];
                            middle <= data2[175:175];
                            right <= data3[175:175];
                        end
                    176:
                        begin
                        left <= data1[176:176];
                            middle <= data2[176:176];
                            right <= data3[176:176];
                        end
                    177:
                        begin
                        left <= data1[177:177];
                            middle <= data2[177:177];
                            right <= data3[177:177];
                        end
                    178:
                        begin
                        left <= data1[178:178];
                            middle <= data2[178:178];
                            right <= data3[178:178];
                        end
                    179:
                        begin
                        left <= data1[179:179];
                            middle <= data2[179:179];
                            right <= data3[179:179];
                        end
                    180:
                        begin
                        left <= data1[180:180];
                            middle <= data2[180:180];
                            right <= data3[180:180];
                        end
                    181:
                        begin
                        left <= data1[181:181];
                            middle <= data2[181:181];
                            right <= data3[181:181];
                        end
                    182:
                        begin
                        left <= data1[182:182];
                            middle <= data2[182:182];
                            right <= data3[182:182];
                        end
                    183:
                        begin
                        left <= data1[183:183];
                            middle <= data2[183:183];
                            right <= data3[183:183];
                        end
                    184:
                        begin
                        left <= data1[184:184];
                            middle <= data2[184:184];
                            right <= data3[184:184];
                        end
                    185:
                        begin
                        left <= data1[185:185];
                            middle <= data2[185:185];
                            right <= data3[185:185];
                        end
                    186:
                        begin
                        left <= data1[186:186];
                            middle <= data2[186:186];
                            right <= data3[186:186];
                        end
                    187:
                        begin
                        left <= data1[187:187];
                            middle <= data2[187:187];
                            right <= data3[187:187];
                        end
                    188:
                        begin
                        left <= data1[188:188];
                            middle <= data2[188:188];
                            right <= data3[188:188];
                        end
                    189:
                        begin
                        left <= data1[189:189];
                            middle <= data2[189:189];
                            right <= data3[189:189];
                        end
                    190:
                        begin
                        left <= data1[190:190];
                            middle <= data2[190:190];
                            right <= data3[190:190];
                        end
                    191:
                        begin
                        left <= data1[191:191];
                            middle <= data2[191:191];
                            right <= data3[191:191];
                        end
                    192:
                        begin
                        left <= data1[192:192];
                            middle <= data2[192:192];
                            right <= data3[192:192];
                        end
                    193:
                        begin
                        left <= data1[193:193];
                            middle <= data2[193:193];
                            right <= data3[193:193];
                        end
                    194:
                        begin
                        left <= data1[194:194];
                            middle <= data2[194:194];
                            right <= data3[194:194];
                        end
                    195:
                        begin
                        left <= data1[195:195];
                            middle <= data2[195:195];
                            right <= data3[195:195];
                        end
                    196:
                        begin
                        left <= data1[196:196];
                            middle <= data2[196:196];
                            right <= data3[196:196];
                        end
                    197:
                        begin
                        left <= data1[197:197];
                            middle <= data2[197:197];
                            right <= data3[197:197];
                        end
                    198:
                        begin
                        left <= data1[198:198];
                            middle <= data2[198:198];
                            right <= data3[198:198];
                        end
                    199:
                        begin
                        left <= data1[199:199];
                            middle <= data2[199:199];
                            right <= data3[199:199];
                        end
                    200:
                        begin
                        left <= data1[200:200];
                            middle <= data2[200:200];
                            right <= data3[200:200];
                        end
                    201:
                        begin
                        left <= data1[201:201];
                            middle <= data2[201:201];
                            right <= data3[201:201];
                        end
                    202:
                        begin
                        left <= data1[202:202];
                            middle <= data2[202:202];
                            right <= data3[202:202];
                        end
                    203:
                        begin
                        left <= data1[203:203];
                            middle <= data2[203:203];
                            right <= data3[203:203];
                        end
                    204:
                        begin
                        left <= data1[204:204];
                            middle <= data2[204:204];
                            right <= data3[204:204];
                        end
                    205:
                        begin
                        left <= data1[205:205];
                            middle <= data2[205:205];
                            right <= data3[205:205];
                        end
                    206:
                        begin
                        left <= data1[206:206];
                            middle <= data2[206:206];
                            right <= data3[206:206];
                        end
                    207:
                        begin
                        left <= data1[207:207];
                            middle <= data2[207:207];
                            right <= data3[207:207];
                        end
                    208:
                        begin
                        left <= data1[208:208];
                            middle <= data2[208:208];
                            right <= data3[208:208];
                        end
                    209:
                        begin
                        left <= data1[209:209];
                            middle <= data2[209:209];
                            right <= data3[209:209];
                        end
                    210:
                        begin
                        left <= data1[210:210];
                            middle <= data2[210:210];
                            right <= data3[210:210];
                        end
                    211:
                        begin
                        left <= data1[211:211];
                            middle <= data2[211:211];
                            right <= data3[211:211];
                        end
                    212:
                        begin
                        left <= data1[212:212];
                            middle <= data2[212:212];
                            right <= data3[212:212];
                        end
                    213:
                        begin
                        left <= data1[213:213];
                            middle <= data2[213:213];
                            right <= data3[213:213];
                        end
                    214:
                        begin
                        left <= data1[214:214];
                            middle <= data2[214:214];
                            right <= data3[214:214];
                        end
                    215:
                        begin
                        left <= data1[215:215];
                            middle <= data2[215:215];
                            right <= data3[215:215];
                        end
                    216:
                        begin
                        left <= data1[216:216];
                            middle <= data2[216:216];
                            right <= data3[216:216];
                        end
                    217:
                        begin
                        left <= data1[217:217];
                            middle <= data2[217:217];
                            right <= data3[217:217];
                        end
                    218:
                        begin
                        left <= data1[218:218];
                            middle <= data2[218:218];
                            right <= data3[218:218];
                        end
                    219:
                        begin
                        left <= data1[219:219];
                            middle <= data2[219:219];
                            right <= data3[219:219];
                        end
                    220:
                        begin
                        left <= data1[220:220];
                            middle <= data2[220:220];
                            right <= data3[220:220];
                        end
                    221:
                        begin
                        left <= data1[221:221];
                            middle <= data2[221:221];
                            right <= data3[221:221];
                        end
                    222:
                        begin
                        left <= data1[222:222];
                            middle <= data2[222:222];
                            right <= data3[222:222];
                        end
                    223:
                        begin
                        left <= data1[223:223];
                            middle <= data2[223:223];
                            right <= data3[223:223];
                        end
                    224:
                        begin
                        left <= data1[224:224];
                            middle <= data2[224:224];
                            right <= data3[224:224];
                        end
                    225:
                        begin
                        left <= data1[225:225];
                            middle <= data2[225:225];
                            right <= data3[225:225];
                        end
                    226:
                        begin
                        left <= data1[226:226];
                            middle <= data2[226:226];
                            right <= data3[226:226];
                        end
                    227:
                        begin
                        left <= data1[227:227];
                            middle <= data2[227:227];
                            right <= data3[227:227];
                        end
                    228:
                        begin
                        left <= data1[228:228];
                            middle <= data2[228:228];
                            right <= data3[228:228];
                        end
                    229:
                        begin
                        left <= data1[229:229];
                            middle <= data2[229:229];
                            right <= data3[229:229];
                        end
                    230:
                        begin
                        left <= data1[230:230];
                            middle <= data2[230:230];
                            right <= data3[230:230];
                        end
                    231:
                        begin
                        left <= data1[231:231];
                            middle <= data2[231:231];
                            right <= data3[231:231];
                        end
                    232:
                        begin
                        left <= data1[232:232];
                            middle <= data2[232:232];
                            right <= data3[232:232];
                        end
                    233:
                        begin
                        left <= data1[233:233];
                            middle <= data2[233:233];
                            right <= data3[233:233];
                        end
                    234:
                        begin
                        left <= data1[234:234];
                            middle <= data2[234:234];
                            right <= data3[234:234];
                        end
                    235:
                        begin
                        left <= data1[235:235];
                            middle <= data2[235:235];
                            right <= data3[235:235];
                        end
                    236:
                        begin
                        left <= data1[236:236];
                            middle <= data2[236:236];
                            right <= data3[236:236];
                        end
                    237:
                        begin
                        left <= data1[237:237];
                            middle <= data2[237:237];
                            right <= data3[237:237];
                        end
                    238:
                        begin
                        left <= data1[238:238];
                            middle <= data2[238:238];
                            right <= data3[238:238];
                        end
                    239:
                        begin
                        left <= data1[239:239];
                            middle <= data2[239:239];
                            right <= data3[239:239];
                        end
                    240:
                        begin
                        left <= data1[240:240];
                            middle <= data2[240:240];
                            right <= data3[240:240];
                        end
                    241:
                        begin
                        left <= data1[241:241];
                            middle <= data2[241:241];
                            right <= data3[241:241];
                        end
                    242:
                        begin
                        left <= data1[242:242];
                            middle <= data2[242:242];
                            right <= data3[242:242];
                        end
                    243:
                        begin
                        left <= data1[243:243];
                            middle <= data2[243:243];
                            right <= data3[243:243];
                        end
                    244:
                        begin
                        left <= data1[244:244];
                            middle <= data2[244:244];
                            right <= data3[244:244];
                        end
                    245:
                        begin
                        left <= data1[245:245];
                            middle <= data2[245:245];
                            right <= data3[245:245];
                        end
                    246:
                        begin
                        left <= data1[246:246];
                            middle <= data2[246:246];
                            right <= data3[246:246];
                        end
                    247:
                        begin
                        left <= data1[247:247];
                            middle <= data2[247:247];
                            right <= data3[247:247];
                        end
                    248:
                        begin
                        left <= data1[248:248];
                            middle <= data2[248:248];
                            right <= data3[248:248];
                        end
                    249:
                        begin
                        left <= data1[249:249];
                            middle <= data2[249:249];
                            right <= data3[249:249];
                        end
                    250:
                        begin
                        left <= data1[250:250];
                            middle <= data2[250:250];
                            right <= data3[250:250];
                        end
                    251:
                        begin
                        left <= data1[251:251];
                            middle <= data2[251:251];
                            right <= data3[251:251];
                        end
                    252:
                        begin
                        left <= data1[252:252];
                            middle <= data2[252:252];
                            right <= data3[252:252];
                        end
                    253:
                        begin
                        left <= data1[253:253];
                            middle <= data2[253:253];
                            right <= data3[253:253];
                        end
                    254:
                        begin
                        left <= data1[254:254];
                            middle <= data2[254:254];
                            right <= data3[254:254];
                        end
                    255:
                        begin
                        left <= data1[255:255];
                            middle <= data2[255:255];
                            right <= data3[255:255];
                        end
                    256:
                        begin
                        left <= data1[256:256];
                            middle <= data2[256:256];
                            right <= data3[256:256];
                        end
                    257:
                        begin
                        left <= data1[257:257];
                            middle <= data2[257:257];
                            right <= data3[257:257];
                        end
                    258:
                        begin
                        left <= data1[258:258];
                            middle <= data2[258:258];
                            right <= data3[258:258];
                        end
                    259:
                        begin
                        left <= data1[259:259];
                            middle <= data2[259:259];
                            right <= data3[259:259];
                        end
                    260:
                        begin
                        left <= data1[260:260];
                            middle <= data2[260:260];
                            right <= data3[260:260];
                        end
                    261:
                        begin
                        left <= data1[261:261];
                            middle <= data2[261:261];
                            right <= data3[261:261];
                        end
                    262:
                        begin
                        left <= data1[262:262];
                            middle <= data2[262:262];
                            right <= data3[262:262];
                        end
                    263:
                        begin
                        left <= data1[263:263];
                            middle <= data2[263:263];
                            right <= data3[263:263];
                        end
                    264:
                        begin
                        left <= data1[264:264];
                            middle <= data2[264:264];
                            right <= data3[264:264];
                        end
                    265:
                        begin
                        left <= data1[265:265];
                            middle <= data2[265:265];
                            right <= data3[265:265];
                        end
                    266:
                        begin
                        left <= data1[266:266];
                            middle <= data2[266:266];
                            right <= data3[266:266];
                        end
                    267:
                        begin
                        left <= data1[267:267];
                            middle <= data2[267:267];
                            right <= data3[267:267];
                        end
                    268:
                        begin
                        left <= data1[268:268];
                            middle <= data2[268:268];
                            right <= data3[268:268];
                        end
                    269:
                        begin
                        left <= data1[269:269];
                            middle <= data2[269:269];
                            right <= data3[269:269];
                        end
                    270:
                        begin
                        left <= data1[270:270];
                            middle <= data2[270:270];
                            right <= data3[270:270];
                        end
                    271:
                        begin
                        left <= data1[271:271];
                            middle <= data2[271:271];
                            right <= data3[271:271];
                        end
                    272:
                        begin
                        left <= data1[272:272];
                            middle <= data2[272:272];
                            right <= data3[272:272];
                        end
                    273:
                        begin
                        left <= data1[273:273];
                            middle <= data2[273:273];
                            right <= data3[273:273];
                        end
                    274:
                        begin
                        left <= data1[274:274];
                            middle <= data2[274:274];
                            right <= data3[274:274];
                        end
                    275:
                        begin
                        left <= data1[275:275];
                            middle <= data2[275:275];
                            right <= data3[275:275];
                        end
                    276:
                        begin
                        left <= data1[276:276];
                            middle <= data2[276:276];
                            right <= data3[276:276];
                        end
                    277:
                        begin
                        left <= data1[277:277];
                            middle <= data2[277:277];
                            right <= data3[277:277];
                        end
                    278:
                        begin
                        left <= data1[278:278];
                            middle <= data2[278:278];
                            right <= data3[278:278];
                        end
                    279:
                        begin
                        left <= data1[279:279];
                            middle <= data2[279:279];
                            right <= data3[279:279];
                        end
                    280:
                        begin
                        left <= data1[280:280];
                            middle <= data2[280:280];
                            right <= data3[280:280];
                        end
                    281:
                        begin
                        left <= data1[281:281];
                            middle <= data2[281:281];
                            right <= data3[281:281];
                        end
                    282:
                        begin
                        left <= data1[282:282];
                            middle <= data2[282:282];
                            right <= data3[282:282];
                        end
                    283:
                        begin
                        left <= data1[283:283];
                            middle <= data2[283:283];
                            right <= data3[283:283];
                        end
                    284:
                        begin
                        left <= data1[284:284];
                            middle <= data2[284:284];
                            right <= data3[284:284];
                        end
                    285:
                        begin
                        left <= data1[285:285];
                            middle <= data2[285:285];
                            right <= data3[285:285];
                        end
                    286:
                        begin
                        left <= data1[286:286];
                            middle <= data2[286:286];
                            right <= data3[286:286];
                        end
                    287:
                        begin
                        left <= data1[287:287];
                            middle <= data2[287:287];
                            right <= data3[287:287];
                        end
                    288:
                        begin
                        left <= data1[288:288];
                            middle <= data2[288:288];
                            right <= data3[288:288];
                        end
                    289:
                        begin
                        left <= data1[289:289];
                            middle <= data2[289:289];
                            right <= data3[289:289];
                        end
                    290:
                        begin
                        left <= data1[290:290];
                            middle <= data2[290:290];
                            right <= data3[290:290];
                        end
                    291:
                        begin
                        left <= data1[291:291];
                            middle <= data2[291:291];
                            right <= data3[291:291];
                        end
                    292:
                        begin
                        left <= data1[292:292];
                            middle <= data2[292:292];
                            right <= data3[292:292];
                        end
                    293:
                        begin
                        left <= data1[293:293];
                            middle <= data2[293:293];
                            right <= data3[293:293];
                        end
                    294:
                        begin
                        left <= data1[294:294];
                            middle <= data2[294:294];
                            right <= data3[294:294];
                        end
                    295:
                        begin
                        left <= data1[295:295];
                            middle <= data2[295:295];
                            right <= data3[295:295];
                        end
                    296:
                        begin
                        left <= data1[296:296];
                            middle <= data2[296:296];
                            right <= data3[296:296];
                        end
                    297:
                        begin
                        left <= data1[297:297];
                            middle <= data2[297:297];
                            right <= data3[297:297];
                        end
                    298:
                        begin
                        left <= data1[298:298];
                            middle <= data2[298:298];
                            right <= data3[298:298];
                        end
                    299:
                        begin
                        left <= data1[299:299];
                            middle <= data2[299:299];
                            right <= data3[299:299];
                        end
                    300:
                        begin
                        left <= data1[300:300];
                            middle <= data2[300:300];
                            right <= data3[300:300];
                        end
                    301:
                        begin
                        left <= data1[301:301];
                            middle <= data2[301:301];
                            right <= data3[301:301];
                        end
                    302:
                        begin
                        left <= data1[302:302];
                            middle <= data2[302:302];
                            right <= data3[302:302];
                        end
                    303:
                        begin
                        left <= data1[303:303];
                            middle <= data2[303:303];
                            right <= data3[303:303];
                        end
                    304:
                        begin
                        left <= data1[304:304];
                            middle <= data2[304:304];
                            right <= data3[304:304];
                        end
                    305:
                        begin
                        left <= data1[305:305];
                            middle <= data2[305:305];
                            right <= data3[305:305];
                        end
                    306:
                        begin
                        left <= data1[306:306];
                            middle <= data2[306:306];
                            right <= data3[306:306];
                        end
                    307:
                        begin
                        left <= data1[307:307];
                            middle <= data2[307:307];
                            right <= data3[307:307];
                        end
                    308:
                        begin
                        left <= data1[308:308];
                            middle <= data2[308:308];
                            right <= data3[308:308];
                        end
                    309:
                        begin
                        left <= data1[309:309];
                            middle <= data2[309:309];
                            right <= data3[309:309];
                        end
                    310:
                        begin
                        left <= data1[310:310];
                            middle <= data2[310:310];
                            right <= data3[310:310];
                        end
                    311:
                        begin
                        left <= data1[311:311];
                            middle <= data2[311:311];
                            right <= data3[311:311];
                        end
                    312:
                        begin
                        left <= data1[312:312];
                            middle <= data2[312:312];
                            right <= data3[312:312];
                        end
                    313:
                        begin
                        left <= data1[313:313];
                            middle <= data2[313:313];
                            right <= data3[313:313];
                        end
                    314:
                        begin
                        left <= data1[314:314];
                            middle <= data2[314:314];
                            right <= data3[314:314];
                        end
                    315:
                        begin
                        left <= data1[315:315];
                            middle <= data2[315:315];
                            right <= data3[315:315];
                        end
                    316:
                        begin
                        left <= data1[316:316];
                            middle <= data2[316:316];
                            right <= data3[316:316];
                        end
                    317:
                        begin
                        left <= data1[317:317];
                            middle <= data2[317:317];
                            right <= data3[317:317];
                        end
                    318:
                        begin
                        left <= data1[318:318];
                            middle <= data2[318:318];
                            right <= data3[318:318];
                        end
                    319:
                        begin
                        left <= data1[319:319];
                            middle <= data2[319:319];
                            right <= data3[319:319];
                        end
                    320:
                        begin
                        left <= data1[320:320];
                            middle <= data2[320:320];
                            right <= data3[320:320];
                        end
                    321:
                        begin
                        left <= data1[321:321];
                            middle <= data2[321:321];
                            right <= data3[321:321];
                        end
                    322:
                        begin
                        left <= data1[322:322];
                            middle <= data2[322:322];
                            right <= data3[322:322];
                        end
                    323:
                        begin
                        left <= data1[323:323];
                            middle <= data2[323:323];
                            right <= data3[323:323];
                        end
                    324:
                        begin
                        left <= data1[324:324];
                            middle <= data2[324:324];
                            right <= data3[324:324];
                        end
                    325:
                        begin
                        left <= data1[325:325];
                            middle <= data2[325:325];
                            right <= data3[325:325];
                        end
                    326:
                        begin
                        left <= data1[326:326];
                            middle <= data2[326:326];
                            right <= data3[326:326];
                        end
                    327:
                        begin
                        left <= data1[327:327];
                            middle <= data2[327:327];
                            right <= data3[327:327];
                        end
                    328:
                        begin
                        left <= data1[328:328];
                            middle <= data2[328:328];
                            right <= data3[328:328];
                        end
                    329:
                        begin
                        left <= data1[329:329];
                            middle <= data2[329:329];
                            right <= data3[329:329];
                        end
                    330:
                        begin
                        left <= data1[330:330];
                            middle <= data2[330:330];
                            right <= data3[330:330];
                        end
                    331:
                        begin
                        left <= data1[331:331];
                            middle <= data2[331:331];
                            right <= data3[331:331];
                        end
                    332:
                        begin
                        left <= data1[332:332];
                            middle <= data2[332:332];
                            right <= data3[332:332];
                        end
                    333:
                        begin
                        left <= data1[333:333];
                            middle <= data2[333:333];
                            right <= data3[333:333];
                        end
                    334:
                        begin
                        left <= data1[334:334];
                            middle <= data2[334:334];
                            right <= data3[334:334];
                        end
                    335:
                        begin
                        left <= data1[335:335];
                            middle <= data2[335:335];
                            right <= data3[335:335];
                        end
                    336:
                        begin
                        left <= data1[336:336];
                            middle <= data2[336:336];
                            right <= data3[336:336];
                        end
                    337:
                        begin
                        left <= data1[337:337];
                            middle <= data2[337:337];
                            right <= data3[337:337];
                        end
                    338:
                        begin
                        left <= data1[338:338];
                            middle <= data2[338:338];
                            right <= data3[338:338];
                        end
                    339:
                        begin
                        left <= data1[339:339];
                            middle <= data2[339:339];
                            right <= data3[339:339];
                        end
                    340:
                        begin
                        left <= data1[340:340];
                            middle <= data2[340:340];
                            right <= data3[340:340];
                        end
                    341:
                        begin
                        left <= data1[341:341];
                            middle <= data2[341:341];
                            right <= data3[341:341];
                        end
                    342:
                        begin
                        left <= data1[342:342];
                            middle <= data2[342:342];
                            right <= data3[342:342];
                        end
                    343:
                        begin
                        left <= data1[343:343];
                            middle <= data2[343:343];
                            right <= data3[343:343];
                        end
                    344:
                        begin
                        left <= data1[344:344];
                            middle <= data2[344:344];
                            right <= data3[344:344];
                        end
                    345:
                        begin
                        left <= data1[345:345];
                            middle <= data2[345:345];
                            right <= data3[345:345];
                        end
                    346:
                        begin
                        left <= data1[346:346];
                            middle <= data2[346:346];
                            right <= data3[346:346];
                        end
                    347:
                        begin
                        left <= data1[347:347];
                            middle <= data2[347:347];
                            right <= data3[347:347];
                        end
                    348:
                        begin
                        left <= data1[348:348];
                            middle <= data2[348:348];
                            right <= data3[348:348];
                        end
                    349:
                        begin
                        left <= data1[349:349];
                            middle <= data2[349:349];
                            right <= data3[349:349];
                        end
                    350:
                        begin
                        left <= data1[350:350];
                            middle <= data2[350:350];
                            right <= data3[350:350];
                        end
                    351:
                        begin
                        left <= data1[351:351];
                            middle <= data2[351:351];
                            right <= data3[351:351];
                        end
                    352:
                        begin
                        left <= data1[352:352];
                            middle <= data2[352:352];
                            right <= data3[352:352];
                        end
                    353:
                        begin
                        left <= data1[353:353];
                            middle <= data2[353:353];
                            right <= data3[353:353];
                        end
                    354:
                        begin
                        left <= data1[354:354];
                            middle <= data2[354:354];
                            right <= data3[354:354];
                        end
                    355:
                        begin
                        left <= data1[355:355];
                            middle <= data2[355:355];
                            right <= data3[355:355];
                        end
                    356:
                        begin
                        left <= data1[356:356];
                            middle <= data2[356:356];
                            right <= data3[356:356];
                        end
                    357:
                        begin
                        left <= data1[357:357];
                            middle <= data2[357:357];
                            right <= data3[357:357];
                        end
                    358:
                        begin
                        left <= data1[358:358];
                            middle <= data2[358:358];
                            right <= data3[358:358];
                        end
                    359:
                        begin
                        left <= data1[359:359];
                            middle <= data2[359:359];
                            right <= data3[359:359];
                        end
                    360:
                        begin
                        left <= data1[360:360];
                            middle <= data2[360:360];
                            right <= data3[360:360];
                        end
                    361:
                        begin
                        left <= data1[361:361];
                            middle <= data2[361:361];
                            right <= data3[361:361];
                        end
                    362:
                        begin
                        left <= data1[362:362];
                            middle <= data2[362:362];
                            right <= data3[362:362];
                        end
                    363:
                        begin
                        left <= data1[363:363];
                            middle <= data2[363:363];
                            right <= data3[363:363];
                        end
                    364:
                        begin
                        left <= data1[364:364];
                            middle <= data2[364:364];
                            right <= data3[364:364];
                        end
                    365:
                        begin
                        left <= data1[365:365];
                            middle <= data2[365:365];
                            right <= data3[365:365];
                        end
                    366:
                        begin
                        left <= data1[366:366];
                            middle <= data2[366:366];
                            right <= data3[366:366];
                        end
                    367:
                        begin
                        left <= data1[367:367];
                            middle <= data2[367:367];
                            right <= data3[367:367];
                        end
                    368:
                        begin
                        left <= data1[368:368];
                            middle <= data2[368:368];
                            right <= data3[368:368];
                        end
                    369:
                        begin
                        left <= data1[369:369];
                            middle <= data2[369:369];
                            right <= data3[369:369];
                        end
                    370:
                        begin
                        left <= data1[370:370];
                            middle <= data2[370:370];
                            right <= data3[370:370];
                        end
                    371:
                        begin
                        left <= data1[371:371];
                            middle <= data2[371:371];
                            right <= data3[371:371];
                        end
                    372:
                        begin
                        left <= data1[372:372];
                            middle <= data2[372:372];
                            right <= data3[372:372];
                        end
                    373:
                        begin
                        left <= data1[373:373];
                            middle <= data2[373:373];
                            right <= data3[373:373];
                        end
                    374:
                        begin
                        left <= data1[374:374];
                            middle <= data2[374:374];
                            right <= data3[374:374];
                        end
                    375:
                        begin
                        left <= data1[375:375];
                            middle <= data2[375:375];
                            right <= data3[375:375];
                        end
                    376:
                        begin
                        left <= data1[376:376];
                            middle <= data2[376:376];
                            right <= data3[376:376];
                        end
                    377:
                        begin
                        left <= data1[377:377];
                            middle <= data2[377:377];
                            right <= data3[377:377];
                        end
                    378:
                        begin
                        left <= data1[378:378];
                            middle <= data2[378:378];
                            right <= data3[378:378];
                        end
                    379:
                        begin
                        left <= data1[379:379];
                            middle <= data2[379:379];
                            right <= data3[379:379];
                        end
                    380:
                        begin
                        left <= data1[380:380];
                            middle <= data2[380:380];
                            right <= data3[380:380];
                        end
                    381:
                        begin
                        left <= data1[381:381];
                            middle <= data2[381:381];
                            right <= data3[381:381];
                        end
                    382:
                        begin
                        left <= data1[382:382];
                            middle <= data2[382:382];
                            right <= data3[382:382];
                        end
                    383:
                        begin
                        left <= data1[383:383];
                            middle <= data2[383:383];
                            right <= data3[383:383];
                        end
                    384:
                        begin
                        left <= data1[384:384];
                            middle <= data2[384:384];
                            right <= data3[384:384];
                        end
                    385:
                        begin
                        left <= data1[385:385];
                            middle <= data2[385:385];
                            right <= data3[385:385];
                        end
                    386:
                        begin
                        left <= data1[386:386];
                            middle <= data2[386:386];
                            right <= data3[386:386];
                        end
                    387:
                        begin
                        left <= data1[387:387];
                            middle <= data2[387:387];
                            right <= data3[387:387];
                        end
                    388:
                        begin
                        left <= data1[388:388];
                            middle <= data2[388:388];
                            right <= data3[388:388];
                        end
                    389:
                        begin
                        left <= data1[389:389];
                            middle <= data2[389:389];
                            right <= data3[389:389];
                        end
                    390:
                        begin
                        left <= data1[390:390];
                            middle <= data2[390:390];
                            right <= data3[390:390];
                        end
                    391:
                        begin
                        left <= data1[391:391];
                            middle <= data2[391:391];
                            right <= data3[391:391];
                        end
                    392:
                        begin
                        left <= data1[392:392];
                            middle <= data2[392:392];
                            right <= data3[392:392];
                        end
                    393:
                        begin
                        left <= data1[393:393];
                            middle <= data2[393:393];
                            right <= data3[393:393];
                        end
                    394:
                        begin
                        left <= data1[394:394];
                            middle <= data2[394:394];
                            right <= data3[394:394];
                        end
                    395:
                        begin
                        left <= data1[395:395];
                            middle <= data2[395:395];
                            right <= data3[395:395];
                        end
                    396:
                        begin
                        left <= data1[396:396];
                            middle <= data2[396:396];
                            right <= data3[396:396];
                        end
                    397:
                        begin
                        left <= data1[397:397];
                            middle <= data2[397:397];
                            right <= data3[397:397];
                        end
                    398:
                        begin
                        left <= data1[398:398];
                            middle <= data2[398:398];
                            right <= data3[398:398];
                        end
                    399:
                        begin
                        left <= data1[399:399];
                            middle <= data2[399:399];
                            right <= data3[399:399];
                        end
                    400:
                        begin
                        left <= data1[400:400];
                            middle <= data2[400:400];
                            right <= data3[400:400];
                        end
                    401:
                        begin
                        left <= data1[401:401];
                            middle <= data2[401:401];
                            right <= data3[401:401];
                        end
                    402:
                        begin
                        left <= data1[402:402];
                            middle <= data2[402:402];
                            right <= data3[402:402];
                        end
                    403:
                        begin
                        left <= data1[403:403];
                            middle <= data2[403:403];
                            right <= data3[403:403];
                        end
                    404:
                        begin
                        left <= data1[404:404];
                            middle <= data2[404:404];
                            right <= data3[404:404];
                        end
                    405:
                        begin
                        left <= data1[405:405];
                            middle <= data2[405:405];
                            right <= data3[405:405];
                        end
                    406:
                        begin
                        left <= data1[406:406];
                            middle <= data2[406:406];
                            right <= data3[406:406];
                        end
                    407:
                        begin
                        left <= data1[407:407];
                            middle <= data2[407:407];
                            right <= data3[407:407];
                        end
                    408:
                        begin
                        left <= data1[408:408];
                            middle <= data2[408:408];
                            right <= data3[408:408];
                        end
                    409:
                        begin
                        left <= data1[409:409];
                            middle <= data2[409:409];
                            right <= data3[409:409];
                        end
                    410:
                        begin
                        left <= data1[410:410];
                            middle <= data2[410:410];
                            right <= data3[410:410];
                        end
                    411:
                        begin
                        left <= data1[411:411];
                            middle <= data2[411:411];
                            right <= data3[411:411];
                        end
                    412:
                        begin
                        left <= data1[412:412];
                            middle <= data2[412:412];
                            right <= data3[412:412];
                        end
                    413:
                        begin
                        left <= data1[413:413];
                            middle <= data2[413:413];
                            right <= data3[413:413];
                        end
                    414:
                        begin
                        left <= data1[414:414];
                            middle <= data2[414:414];
                            right <= data3[414:414];
                        end
                    415:
                        begin
                        left <= data1[415:415];
                            middle <= data2[415:415];
                            right <= data3[415:415];
                        end
                    416:
                        begin
                        left <= data1[416:416];
                            middle <= data2[416:416];
                            right <= data3[416:416];
                        end
                    417:
                        begin
                        left <= data1[417:417];
                            middle <= data2[417:417];
                            right <= data3[417:417];
                        end
                    418:
                        begin
                        left <= data1[418:418];
                            middle <= data2[418:418];
                            right <= data3[418:418];
                        end
                    419:
                        begin
                        left <= data1[419:419];
                            middle <= data2[419:419];
                            right <= data3[419:419];
                        end
                    420:
                        begin
                        left <= data1[420:420];
                            middle <= data2[420:420];
                            right <= data3[420:420];
                        end
                    421:
                        begin
                        left <= data1[421:421];
                            middle <= data2[421:421];
                            right <= data3[421:421];
                        end
                    422:
                        begin
                        left <= data1[422:422];
                            middle <= data2[422:422];
                            right <= data3[422:422];
                        end
                    423:
                        begin
                        left <= data1[423:423];
                            middle <= data2[423:423];
                            right <= data3[423:423];
                        end
                    424:
                        begin
                        left <= data1[424:424];
                            middle <= data2[424:424];
                            right <= data3[424:424];
                        end
                    425:
                        begin
                        left <= data1[425:425];
                            middle <= data2[425:425];
                            right <= data3[425:425];
                        end
                    426:
                        begin
                        left <= data1[426:426];
                            middle <= data2[426:426];
                            right <= data3[426:426];
                        end
                    427:
                        begin
                        left <= data1[427:427];
                            middle <= data2[427:427];
                            right <= data3[427:427];
                        end
                    428:
                        begin
                        left <= data1[428:428];
                            middle <= data2[428:428];
                            right <= data3[428:428];
                        end
                    429:
                        begin
                        left <= data1[429:429];
                            middle <= data2[429:429];
                            right <= data3[429:429];
                        end
                    430:
                        begin
                        left <= data1[430:430];
                            middle <= data2[430:430];
                            right <= data3[430:430];
                        end
                    431:
                        begin
                        left <= data1[431:431];
                            middle <= data2[431:431];
                            right <= data3[431:431];
                        end
                    432:
                        begin
                        left <= data1[432:432];
                            middle <= data2[432:432];
                            right <= data3[432:432];
                        end
                    433:
                        begin
                        left <= data1[433:433];
                            middle <= data2[433:433];
                            right <= data3[433:433];
                        end
                    434:
                        begin
                        left <= data1[434:434];
                            middle <= data2[434:434];
                            right <= data3[434:434];
                        end
                    435:
                        begin
                        left <= data1[435:435];
                            middle <= data2[435:435];
                            right <= data3[435:435];
                        end
                    436:
                        begin
                        left <= data1[436:436];
                            middle <= data2[436:436];
                            right <= data3[436:436];
                        end
                    437:
                        begin
                        left <= data1[437:437];
                            middle <= data2[437:437];
                            right <= data3[437:437];
                        end
                    438:
                        begin
                        left <= data1[438:438];
                            middle <= data2[438:438];
                            right <= data3[438:438];
                        end
                    439:
                        begin
                        left <= data1[439:439];
                            middle <= data2[439:439];
                            right <= data3[439:439];
                        end
                    440:
                        begin
                        left <= data1[440:440];
                            middle <= data2[440:440];
                            right <= data3[440:440];
                        end
                    441:
                        begin
                        left <= data1[441:441];
                            middle <= data2[441:441];
                            right <= data3[441:441];
                        end
                    442:
                        begin
                        left <= data1[442:442];
                            middle <= data2[442:442];
                            right <= data3[442:442];
                        end
                    443:
                        begin
                        left <= data1[443:443];
                            middle <= data2[443:443];
                            right <= data3[443:443];
                        end
                    444:
                        begin
                        left <= data1[444:444];
                            middle <= data2[444:444];
                            right <= data3[444:444];
                        end
                    445:
                        begin
                        left <= data1[445:445];
                            middle <= data2[445:445];
                            right <= data3[445:445];
                        end
                    446:
                        begin
                        left <= data1[446:446];
                            middle <= data2[446:446];
                            right <= data3[446:446];
                        end
                    447:
                        begin
                        left <= data1[447:447];
                            middle <= data2[447:447];
                            right <= data3[447:447];
                        end
                    448:
                        begin
                        left <= data1[448:448];
                            middle <= data2[448:448];
                            right <= data3[448:448];
                        end
                    449:
                        begin
                        left <= data1[449:449];
                            middle <= data2[449:449];
                            right <= data3[449:449];
                        end
                    450:
                        begin
                        left <= data1[450:450];
                            middle <= data2[450:450];
                            right <= data3[450:450];
                        end
                    451:
                        begin
                        left <= data1[451:451];
                            middle <= data2[451:451];
                            right <= data3[451:451];
                        end
                    452:
                        begin
                        left <= data1[452:452];
                            middle <= data2[452:452];
                            right <= data3[452:452];
                        end
                    453:
                        begin
                        left <= data1[453:453];
                            middle <= data2[453:453];
                            right <= data3[453:453];
                        end
                    454:
                        begin
                        left <= data1[454:454];
                            middle <= data2[454:454];
                            right <= data3[454:454];
                        end
                    455:
                        begin
                        left <= data1[455:455];
                            middle <= data2[455:455];
                            right <= data3[455:455];
                        end
                    456:
                        begin
                        left <= data1[456:456];
                            middle <= data2[456:456];
                            right <= data3[456:456];
                        end
                    457:
                        begin
                        left <= data1[457:457];
                            middle <= data2[457:457];
                            right <= data3[457:457];
                        end
                    458:
                        begin
                        left <= data1[458:458];
                            middle <= data2[458:458];
                            right <= data3[458:458];
                        end
                    459:
                        begin
                        left <= data1[459:459];
                            middle <= data2[459:459];
                            right <= data3[459:459];
                        end
                    460:
                        begin
                        left <= data1[460:460];
                            middle <= data2[460:460];
                            right <= data3[460:460];
                        end
                    461:
                        begin
                        left <= data1[461:461];
                            middle <= data2[461:461];
                            right <= data3[461:461];
                        end
                    462:
                        begin
                        left <= data1[462:462];
                            middle <= data2[462:462];
                            right <= data3[462:462];
                        end
                    463:
                        begin
                        left <= data1[463:463];
                            middle <= data2[463:463];
                            right <= data3[463:463];
                        end
                    464:
                        begin
                        left <= data1[464:464];
                            middle <= data2[464:464];
                            right <= data3[464:464];
                        end
                    465:
                        begin
                        left <= data1[465:465];
                            middle <= data2[465:465];
                            right <= data3[465:465];
                        end
                    466:
                        begin
                        left <= data1[466:466];
                            middle <= data2[466:466];
                            right <= data3[466:466];
                        end
                    467:
                        begin
                        left <= data1[467:467];
                            middle <= data2[467:467];
                            right <= data3[467:467];
                        end
                    468:
                        begin
                        left <= data1[468:468];
                            middle <= data2[468:468];
                            right <= data3[468:468];
                        end
                    469:
                        begin
                        left <= data1[469:469];
                            middle <= data2[469:469];
                            right <= data3[469:469];
                        end
                    470:
                        begin
                        left <= data1[470:470];
                            middle <= data2[470:470];
                            right <= data3[470:470];
                        end
                    471:
                        begin
                        left <= data1[471:471];
                            middle <= data2[471:471];
                            right <= data3[471:471];
                        end
                    472:
                        begin
                        left <= data1[472:472];
                            middle <= data2[472:472];
                            right <= data3[472:472];
                        end
                    473:
                        begin
                        left <= data1[473:473];
                            middle <= data2[473:473];
                            right <= data3[473:473];
                        end
                    474:
                        begin
                        left <= data1[474:474];
                            middle <= data2[474:474];
                            right <= data3[474:474];
                        end
                    475:
                        begin
                        left <= data1[475:475];
                            middle <= data2[475:475];
                            right <= data3[475:475];
                        end
                    476:
                        begin
                        left <= data1[476:476];
                            middle <= data2[476:476];
                            right <= data3[476:476];
                        end
                    477:
                        begin
                        left <= data1[477:477];
                            middle <= data2[477:477];
                            right <= data3[477:477];
                        end
                    478:
                        begin
                        left <= data1[478:478];
                            middle <= data2[478:478];
                            right <= data3[478:478];
                        end
                    479:
                        begin
                        left <= data1[479:479];
                            middle <= data2[479:479];
                            right <= data3[479:479];
                        end
                    480:
                        begin
                        left <= data1[480:480];
                            middle <= data2[480:480];
                            right <= data3[480:480];
                        end
                    481:
                        begin
                        left <= data1[481:481];
                            middle <= data2[481:481];
                            right <= data3[481:481];
                        end
                    482:
                        begin
                        left <= data1[482:482];
                            middle <= data2[482:482];
                            right <= data3[482:482];
                        end
                    483:
                        begin
                        left <= data1[483:483];
                            middle <= data2[483:483];
                            right <= data3[483:483];
                        end
                    484:
                        begin
                        left <= data1[484:484];
                            middle <= data2[484:484];
                            right <= data3[484:484];
                        end
                    485:
                        begin
                        left <= data1[485:485];
                            middle <= data2[485:485];
                            right <= data3[485:485];
                        end
                    486:
                        begin
                        left <= data1[486:486];
                            middle <= data2[486:486];
                            right <= data3[486:486];
                        end
                    487:
                        begin
                        left <= data1[487:487];
                            middle <= data2[487:487];
                            right <= data3[487:487];
                        end
                    488:
                        begin
                        left <= data1[488:488];
                            middle <= data2[488:488];
                            right <= data3[488:488];
                        end
                    489:
                        begin
                        left <= data1[489:489];
                            middle <= data2[489:489];
                            right <= data3[489:489];
                        end
                    490:
                        begin
                        left <= data1[490:490];
                            middle <= data2[490:490];
                            right <= data3[490:490];
                        end
                    491:
                        begin
                        left <= data1[491:491];
                            middle <= data2[491:491];
                            right <= data3[491:491];
                        end
                    492:
                        begin
                        left <= data1[492:492];
                            middle <= data2[492:492];
                            right <= data3[492:492];
                        end
                    493:
                        begin
                        left <= data1[493:493];
                            middle <= data2[493:493];
                            right <= data3[493:493];
                        end
                    494:
                        begin
                        left <= data1[494:494];
                            middle <= data2[494:494];
                            right <= data3[494:494];
                        end
                    495:
                        begin
                        left <= data1[495:495];
                            middle <= data2[495:495];
                            right <= data3[495:495];
                        end
                    496:
                        begin
                        left <= data1[496:496];
                            middle <= data2[496:496];
                            right <= data3[496:496];
                        end
                    497:
                        begin
                        left <= data1[497:497];
                            middle <= data2[497:497];
                            right <= data3[497:497];
                        end
                    498:
                        begin
                        left <= data1[498:498];
                            middle <= data2[498:498];
                            right <= data3[498:498];
                        end
                    499:
                        begin
                        left <= data1[499:499];
                            middle <= data2[499:499];
                            right <= data3[499:499];
                        end
                    500:
                        begin
                        left <= data1[500:500];
                            middle <= data2[500:500];
                            right <= data3[500:500];
                        end
                    501:
                        begin
                        left <= data1[501:501];
                            middle <= data2[501:501];
                            right <= data3[501:501];
                        end
                    502:
                        begin
                        left <= data1[502:502];
                            middle <= data2[502:502];
                            right <= data3[502:502];
                        end
                    503:
                        begin
                        left <= data1[503:503];
                            middle <= data2[503:503];
                            right <= data3[503:503];
                        end
                    504:
                        begin
                        left <= data1[504:504];
                            middle <= data2[504:504];
                            right <= data3[504:504];
                        end
                    505:
                        begin
                        left <= data1[505:505];
                            middle <= data2[505:505];
                            right <= data3[505:505];
                        end
                    506:
                        begin
                        left <= data1[506:506];
                            middle <= data2[506:506];
                            right <= data3[506:506];
                        end
                    507:
                        begin
                        left <= data1[507:507];
                            middle <= data2[507:507];
                            right <= data3[507:507];
                        end
                    508:
                        begin
                        left <= data1[508:508];
                            middle <= data2[508:508];
                            right <= data3[508:508];
                        end
                    509:
                        begin
                        left <= data1[509:509];
                            middle <= data2[509:509];
                            right <= data3[509:509];
                        end
                    510:
                        begin
                        left <= data1[510:510];
                            middle <= data2[510:510];
                            right <= data3[510:510];
                        end
                    511:
                        begin
                        left <= data1[511:511];
                            middle <= data2[511:511];
                            right <= data3[511:511];
                        end
                    512:
                        begin
                        left <= data1[512:512];
                            middle <= data2[512:512];
                            right <= data3[512:512];
                        end
                    513:
                        begin
                        left <= data1[513:513];
                            middle <= data2[513:513];
                            right <= data3[513:513];
                        end
                    514:
                        begin
                        left <= data1[514:514];
                            middle <= data2[514:514];
                            right <= data3[514:514];
                        end
                    515:
                        begin
                        left <= data1[515:515];
                            middle <= data2[515:515];
                            right <= data3[515:515];
                        end
                    516:
                        begin
                        left <= data1[516:516];
                            middle <= data2[516:516];
                            right <= data3[516:516];
                        end
                    517:
                        begin
                        left <= data1[517:517];
                            middle <= data2[517:517];
                            right <= data3[517:517];
                        end
                    518:
                        begin
                        left <= data1[518:518];
                            middle <= data2[518:518];
                            right <= data3[518:518];
                        end
                    519:
                        begin
                        left <= data1[519:519];
                            middle <= data2[519:519];
                            right <= data3[519:519];
                        end
                    520:
                        begin
                        left <= data1[520:520];
                            middle <= data2[520:520];
                            right <= data3[520:520];
                        end
                    521:
                        begin
                        left <= data1[521:521];
                            middle <= data2[521:521];
                            right <= data3[521:521];
                        end
                    522:
                        begin
                        left <= data1[522:522];
                            middle <= data2[522:522];
                            right <= data3[522:522];
                        end
                    523:
                        begin
                        left <= data1[523:523];
                            middle <= data2[523:523];
                            right <= data3[523:523];
                        end
                    524:
                        begin
                        left <= data1[524:524];
                            middle <= data2[524:524];
                            right <= data3[524:524];
                        end
                    525:
                        begin
                        left <= data1[525:525];
                            middle <= data2[525:525];
                            right <= data3[525:525];
                        end
                    526:
                        begin
                        left <= data1[526:526];
                            middle <= data2[526:526];
                            right <= data3[526:526];
                        end
                    527:
                        begin
                        left <= data1[527:527];
                            middle <= data2[527:527];
                            right <= data3[527:527];
                        end
                    528:
                        begin
                        left <= data1[528:528];
                            middle <= data2[528:528];
                            right <= data3[528:528];
                        end
                    529:
                        begin
                        left <= data1[529:529];
                            middle <= data2[529:529];
                            right <= data3[529:529];
                        end
                    530:
                        begin
                        left <= data1[530:530];
                            middle <= data2[530:530];
                            right <= data3[530:530];
                        end
                    531:
                        begin
                        left <= data1[531:531];
                            middle <= data2[531:531];
                            right <= data3[531:531];
                        end
                    532:
                        begin
                        left <= data1[532:532];
                            middle <= data2[532:532];
                            right <= data3[532:532];
                        end
                    533:
                        begin
                        left <= data1[533:533];
                            middle <= data2[533:533];
                            right <= data3[533:533];
                        end
                    534:
                        begin
                        left <= data1[534:534];
                            middle <= data2[534:534];
                            right <= data3[534:534];
                        end
                    535:
                        begin
                        left <= data1[535:535];
                            middle <= data2[535:535];
                            right <= data3[535:535];
                        end
                    536:
                        begin
                        left <= data1[536:536];
                            middle <= data2[536:536];
                            right <= data3[536:536];
                        end
                    537:
                        begin
                        left <= data1[537:537];
                            middle <= data2[537:537];
                            right <= data3[537:537];
                        end
                    538:
                        begin
                        left <= data1[538:538];
                            middle <= data2[538:538];
                            right <= data3[538:538];
                        end
                    539:
                        begin
                        left <= data1[539:539];
                            middle <= data2[539:539];
                            right <= data3[539:539];
                        end
                    540:
                        begin
                        left <= data1[540:540];
                            middle <= data2[540:540];
                            right <= data3[540:540];
                        end
                    541:
                        begin
                        left <= data1[541:541];
                            middle <= data2[541:541];
                            right <= data3[541:541];
                        end
                    542:
                        begin
                        left <= data1[542:542];
                            middle <= data2[542:542];
                            right <= data3[542:542];
                        end
                    543:
                        begin
                        left <= data1[543:543];
                            middle <= data2[543:543];
                            right <= data3[543:543];
                        end
                    544:
                        begin
                        left <= data1[544:544];
                            middle <= data2[544:544];
                            right <= data3[544:544];
                        end
                    545:
                        begin
                        left <= data1[545:545];
                            middle <= data2[545:545];
                            right <= data3[545:545];
                        end
                    546:
                        begin
                        left <= data1[546:546];
                            middle <= data2[546:546];
                            right <= data3[546:546];
                        end
                    547:
                        begin
                        left <= data1[547:547];
                            middle <= data2[547:547];
                            right <= data3[547:547];
                        end
                    548:
                        begin
                        left <= data1[548:548];
                            middle <= data2[548:548];
                            right <= data3[548:548];
                        end
                    549:
                        begin
                        left <= data1[549:549];
                            middle <= data2[549:549];
                            right <= data3[549:549];
                        end
                    550:
                        begin
                        left <= data1[550:550];
                            middle <= data2[550:550];
                            right <= data3[550:550];
                        end
                    551:
                        begin
                        left <= data1[551:551];
                            middle <= data2[551:551];
                            right <= data3[551:551];
                        end
                    552:
                        begin
                        left <= data1[552:552];
                            middle <= data2[552:552];
                            right <= data3[552:552];
                        end
                    553:
                        begin
                        left <= data1[553:553];
                            middle <= data2[553:553];
                            right <= data3[553:553];
                        end
                    554:
                        begin
                        left <= data1[554:554];
                            middle <= data2[554:554];
                            right <= data3[554:554];
                        end
                    555:
                        begin
                        left <= data1[555:555];
                            middle <= data2[555:555];
                            right <= data3[555:555];
                        end
                    556:
                        begin
                        left <= data1[556:556];
                            middle <= data2[556:556];
                            right <= data3[556:556];
                        end
                    557:
                        begin
                        left <= data1[557:557];
                            middle <= data2[557:557];
                            right <= data3[557:557];
                        end
                    558:
                        begin
                        left <= data1[558:558];
                            middle <= data2[558:558];
                            right <= data3[558:558];
                        end
                    559:
                        begin
                        left <= data1[559:559];
                            middle <= data2[559:559];
                            right <= data3[559:559];
                        end
                    560:
                        begin
                        left <= data1[560:560];
                            middle <= data2[560:560];
                            right <= data3[560:560];
                        end
                    561:
                        begin
                        left <= data1[561:561];
                            middle <= data2[561:561];
                            right <= data3[561:561];
                        end
                    562:
                        begin
                        left <= data1[562:562];
                            middle <= data2[562:562];
                            right <= data3[562:562];
                        end
                    563:
                        begin
                        left <= data1[563:563];
                            middle <= data2[563:563];
                            right <= data3[563:563];
                        end
                    564:
                        begin
                        left <= data1[564:564];
                            middle <= data2[564:564];
                            right <= data3[564:564];
                        end
                    565:
                        begin
                        left <= data1[565:565];
                            middle <= data2[565:565];
                            right <= data3[565:565];
                        end
                    566:
                        begin
                        left <= data1[566:566];
                            middle <= data2[566:566];
                            right <= data3[566:566];
                        end
                    567:
                        begin
                        left <= data1[567:567];
                            middle <= data2[567:567];
                            right <= data3[567:567];
                        end
                    568:
                        begin
                        left <= data1[568:568];
                            middle <= data2[568:568];
                            right <= data3[568:568];
                        end
                    569:
                        begin
                        left <= data1[569:569];
                            middle <= data2[569:569];
                            right <= data3[569:569];
                        end
                    570:
                        begin
                        left <= data1[570:570];
                            middle <= data2[570:570];
                            right <= data3[570:570];
                        end
                    571:
                        begin
                        left <= data1[571:571];
                            middle <= data2[571:571];
                            right <= data3[571:571];
                        end
                    572:
                        begin
                        left <= data1[572:572];
                            middle <= data2[572:572];
                            right <= data3[572:572];
                        end
                    573:
                        begin
                        left <= data1[573:573];
                            middle <= data2[573:573];
                            right <= data3[573:573];
                        end
                    574:
                        begin
                        left <= data1[574:574];
                            middle <= data2[574:574];
                            right <= data3[574:574];
                        end
                    575:
                        begin
                        left <= data1[575:575];
                            middle <= data2[575:575];
                            right <= data3[575:575];
                        end
                    576:
                        begin
                        left <= data1[576:576];
                            middle <= data2[576:576];
                            right <= data3[576:576];
                        end
                    577:
                        begin
                        left <= data1[577:577];
                            middle <= data2[577:577];
                            right <= data3[577:577];
                        end
                    578:
                        begin
                        left <= data1[578:578];
                            middle <= data2[578:578];
                            right <= data3[578:578];
                        end
                    579:
                        begin
                        left <= data1[579:579];
                            middle <= data2[579:579];
                            right <= data3[579:579];
                        end
                    580:
                        begin
                        left <= data1[580:580];
                            middle <= data2[580:580];
                            right <= data3[580:580];
                        end
                    581:
                        begin
                        left <= data1[581:581];
                            middle <= data2[581:581];
                            right <= data3[581:581];
                        end
                    582:
                        begin
                        left <= data1[582:582];
                            middle <= data2[582:582];
                            right <= data3[582:582];
                        end
                    583:
                        begin
                        left <= data1[583:583];
                            middle <= data2[583:583];
                            right <= data3[583:583];
                        end
                    584:
                        begin
                        left <= data1[584:584];
                            middle <= data2[584:584];
                            right <= data3[584:584];
                        end
                    585:
                        begin
                        left <= data1[585:585];
                            middle <= data2[585:585];
                            right <= data3[585:585];
                        end
                    586:
                        begin
                        left <= data1[586:586];
                            middle <= data2[586:586];
                            right <= data3[586:586];
                        end
                    587:
                        begin
                        left <= data1[587:587];
                            middle <= data2[587:587];
                            right <= data3[587:587];
                        end
                    588:
                        begin
                        left <= data1[588:588];
                            middle <= data2[588:588];
                            right <= data3[588:588];
                        end
                    589:
                        begin
                        left <= data1[589:589];
                            middle <= data2[589:589];
                            right <= data3[589:589];
                        end
                    590:
                        begin
                        left <= data1[590:590];
                            middle <= data2[590:590];
                            right <= data3[590:590];
                        end
                    591:
                        begin
                        left <= data1[591:591];
                            middle <= data2[591:591];
                            right <= data3[591:591];
                        end
                    592:
                        begin
                        left <= data1[592:592];
                            middle <= data2[592:592];
                            right <= data3[592:592];
                        end
                    593:
                        begin
                        left <= data1[593:593];
                            middle <= data2[593:593];
                            right <= data3[593:593];
                        end
                    594:
                        begin
                        left <= data1[594:594];
                            middle <= data2[594:594];
                            right <= data3[594:594];
                        end
                    595:
                        begin
                        left <= data1[595:595];
                            middle <= data2[595:595];
                            right <= data3[595:595];
                        end
                    596:
                        begin
                        left <= data1[596:596];
                            middle <= data2[596:596];
                            right <= data3[596:596];
                        end
                    597:
                        begin
                        left <= data1[597:597];
                            middle <= data2[597:597];
                            right <= data3[597:597];
                        end
                    598:
                        begin
                        left <= data1[598:598];
                            middle <= data2[598:598];
                            right <= data3[598:598];
                        end
                    599:
                        begin
                        left <= data1[599:599];
                            middle <= data2[599:599];
                            right <= data3[599:599];
                        end
                    600:
                        begin
                        left <= data1[600:600];
                            middle <= data2[600:600];
                            right <= data3[600:600];
                        end
                    601:
                        begin
                        left <= data1[601:601];
                            middle <= data2[601:601];
                            right <= data3[601:601];
                        end
                    602:
                        begin
                        left <= data1[602:602];
                            middle <= data2[602:602];
                            right <= data3[602:602];
                        end
                    603:
                        begin
                        left <= data1[603:603];
                            middle <= data2[603:603];
                            right <= data3[603:603];
                        end
                    604:
                        begin
                        left <= data1[604:604];
                            middle <= data2[604:604];
                            right <= data3[604:604];
                        end
                    605:
                        begin
                        left <= data1[605:605];
                            middle <= data2[605:605];
                            right <= data3[605:605];
                        end
                    606:
                        begin
                        left <= data1[606:606];
                            middle <= data2[606:606];
                            right <= data3[606:606];
                        end
                    607:
                        begin
                        left <= data1[607:607];
                            middle <= data2[607:607];
                            right <= data3[607:607];
                        end
                    608:
                        begin
                        left <= data1[608:608];
                            middle <= data2[608:608];
                            right <= data3[608:608];
                        end
                    609:
                        begin
                        left <= data1[609:609];
                            middle <= data2[609:609];
                            right <= data3[609:609];
                        end
                    610:
                        begin
                        left <= data1[610:610];
                            middle <= data2[610:610];
                            right <= data3[610:610];
                        end
                    611:
                        begin
                        left <= data1[611:611];
                            middle <= data2[611:611];
                            right <= data3[611:611];
                        end
                    612:
                        begin
                        left <= data1[612:612];
                            middle <= data2[612:612];
                            right <= data3[612:612];
                        end
                    613:
                        begin
                        left <= data1[613:613];
                            middle <= data2[613:613];
                            right <= data3[613:613];
                        end
                    614:
                        begin
                        left <= data1[614:614];
                            middle <= data2[614:614];
                            right <= data3[614:614];
                        end
                    615:
                        begin
                        left <= data1[615:615];
                            middle <= data2[615:615];
                            right <= data3[615:615];
                        end
                    616:
                        begin
                        left <= data1[616:616];
                            middle <= data2[616:616];
                            right <= data3[616:616];
                        end
                    617:
                        begin
                        left <= data1[617:617];
                            middle <= data2[617:617];
                            right <= data3[617:617];
                        end
                    618:
                        begin
                        left <= data1[618:618];
                            middle <= data2[618:618];
                            right <= data3[618:618];
                        end
                    619:
                        begin
                        left <= data1[619:619];
                            middle <= data2[619:619];
                            right <= data3[619:619];
                        end
                    620:
                        begin
                        left <= data1[620:620];
                            middle <= data2[620:620];
                            right <= data3[620:620];
                        end
                    621:
                        begin
                        left <= data1[621:621];
                            middle <= data2[621:621];
                            right <= data3[621:621];
                        end
                    622:
                        begin
                        left <= data1[622:622];
                            middle <= data2[622:622];
                            right <= data3[622:622];
                        end
                    623:
                        begin
                        left <= data1[623:623];
                            middle <= data2[623:623];
                            right <= data3[623:623];
                        end
                    624:
                        begin
                        left <= data1[624:624];
                            middle <= data2[624:624];
                            right <= data3[624:624];
                        end
                    625:
                        begin
                        left <= data1[625:625];
                            middle <= data2[625:625];
                            right <= data3[625:625];
                        end
                    626:
                        begin
                        left <= data1[626:626];
                            middle <= data2[626:626];
                            right <= data3[626:626];
                        end
                    627:
                        begin
                        left <= data1[627:627];
                            middle <= data2[627:627];
                            right <= data3[627:627];
                        end
                    628:
                        begin
                        left <= data1[628:628];
                            middle <= data2[628:628];
                            right <= data3[628:628];
                        end
                    629:
                        begin
                        left <= data1[629:629];
                            middle <= data2[629:629];
                            right <= data3[629:629];
                        end
                    630:
                        begin
                        left <= data1[630:630];
                            middle <= data2[630:630];
                            right <= data3[630:630];
                        end
                    631:
                        begin
                        left <= data1[631:631];
                            middle <= data2[631:631];
                            right <= data3[631:631];
                        end
                    632:
                        begin
                        left <= data1[632:632];
                            middle <= data2[632:632];
                            right <= data3[632:632];
                        end
                    633:
                        begin
                        left <= data1[633:633];
                            middle <= data2[633:633];
                            right <= data3[633:633];
                        end
                    634:
                        begin
                        left <= data1[634:634];
                            middle <= data2[634:634];
                            right <= data3[634:634];
                        end
                    635:
                        begin
                        left <= data1[635:635];
                            middle <= data2[635:635];
                            right <= data3[635:635];
                        end
                    636:
                        begin
                        left <= data1[636:636];
                            middle <= data2[636:636];
                            right <= data3[636:636];
                        end
                    637:
                        begin
                        left <= data1[637:637];
                            middle <= data2[637:637];
                            right <= data3[637:637];
                        end
                    638:
                        begin
                        left <= data1[638:638];
                            middle <= data2[638:638];
                            right <= data3[638:638];
                        end
                    639:
                        begin
                        left <= data1[639:639];
                            middle <= data2[639:639];
                            right <= data3[639:639];
                        end
                    640:
                        begin
                        left <= data1[640:640];
                            middle <= data2[640:640];
                            right <= data3[640:640];
                        end
                    641:
                        begin
                        left <= data1[641:641];
                            middle <= data2[641:641];
                            right <= data3[641:641];
                        end
                    642:
                        begin
                        left <= data1[642:642];
                            middle <= data2[642:642];
                            right <= data3[642:642];
                        end
                    643:
                        begin
                        left <= data1[643:643];
                            middle <= data2[643:643];
                            right <= data3[643:643];
                        end
                    644:
                        begin
                        left <= data1[644:644];
                            middle <= data2[644:644];
                            right <= data3[644:644];
                        end
                    645:
                        begin
                        left <= data1[645:645];
                            middle <= data2[645:645];
                            right <= data3[645:645];
                        end
                    646:
                        begin
                        left <= data1[646:646];
                            middle <= data2[646:646];
                            right <= data3[646:646];
                        end
                    647:
                        begin
                        left <= data1[647:647];
                            middle <= data2[647:647];
                            right <= data3[647:647];
                        end
                    648:
                        begin
                        left <= data1[648:648];
                            middle <= data2[648:648];
                            right <= data3[648:648];
                        end
                    649:
                        begin
                        left <= data1[649:649];
                            middle <= data2[649:649];
                            right <= data3[649:649];
                        end
                    650:
                        begin
                        left <= data1[650:650];
                            middle <= data2[650:650];
                            right <= data3[650:650];
                        end
                    651:
                        begin
                        left <= data1[651:651];
                            middle <= data2[651:651];
                            right <= data3[651:651];
                        end
                    652:
                        begin
                        left <= data1[652:652];
                            middle <= data2[652:652];
                            right <= data3[652:652];
                        end
                    653:
                        begin
                        left <= data1[653:653];
                            middle <= data2[653:653];
                            right <= data3[653:653];
                        end
                    654:
                        begin
                        left <= data1[654:654];
                            middle <= data2[654:654];
                            right <= data3[654:654];
                        end
                    655:
                        begin
                        left <= data1[655:655];
                            middle <= data2[655:655];
                            right <= data3[655:655];
                        end
                    656:
                        begin
                        left <= data1[656:656];
                            middle <= data2[656:656];
                            right <= data3[656:656];
                        end
                    657:
                        begin
                        left <= data1[657:657];
                            middle <= data2[657:657];
                            right <= data3[657:657];
                        end
                    658:
                        begin
                        left <= data1[658:658];
                            middle <= data2[658:658];
                            right <= data3[658:658];
                        end
                    659:
                        begin
                        left <= data1[659:659];
                            middle <= data2[659:659];
                            right <= data3[659:659];
                        end
                    660:
                        begin
                        left <= data1[660:660];
                            middle <= data2[660:660];
                            right <= data3[660:660];
                        end
                    661:
                        begin
                        left <= data1[661:661];
                            middle <= data2[661:661];
                            right <= data3[661:661];
                        end
                    662:
                        begin
                        left <= data1[662:662];
                            middle <= data2[662:662];
                            right <= data3[662:662];
                        end
                    663:
                        begin
                        left <= data1[663:663];
                            middle <= data2[663:663];
                            right <= data3[663:663];
                        end
                    664:
                        begin
                        left <= data1[664:664];
                            middle <= data2[664:664];
                            right <= data3[664:664];
                        end
                    665:
                        begin
                        left <= data1[665:665];
                            middle <= data2[665:665];
                            right <= data3[665:665];
                        end
                    666:
                        begin
                        left <= data1[666:666];
                            middle <= data2[666:666];
                            right <= data3[666:666];
                        end
                    667:
                        begin
                        left <= data1[667:667];
                            middle <= data2[667:667];
                            right <= data3[667:667];
                        end
                    668:
                        begin
                        left <= data1[668:668];
                            middle <= data2[668:668];
                            right <= data3[668:668];
                        end
                    669:
                        begin
                        left <= data1[669:669];
                            middle <= data2[669:669];
                            right <= data3[669:669];
                        end
                    670:
                        begin
                        left <= data1[670:670];
                            middle <= data2[670:670];
                            right <= data3[670:670];
                        end
                    671:
                        begin
                        left <= data1[671:671];
                            middle <= data2[671:671];
                            right <= data3[671:671];
                        end
                    672:
                        begin
                        left <= data1[672:672];
                            middle <= data2[672:672];
                            right <= data3[672:672];
                        end
                    673:
                        begin
                        left <= data1[673:673];
                            middle <= data2[673:673];
                            right <= data3[673:673];
                        end
                    674:
                        begin
                        left <= data1[674:674];
                            middle <= data2[674:674];
                            right <= data3[674:674];
                        end
                    675:
                        begin
                        left <= data1[675:675];
                            middle <= data2[675:675];
                            right <= data3[675:675];
                        end
                    676:
                        begin
                        left <= data1[676:676];
                            middle <= data2[676:676];
                            right <= data3[676:676];
                        end
                    677:
                        begin
                        left <= data1[677:677];
                            middle <= data2[677:677];
                            right <= data3[677:677];
                        end
                    678:
                        begin
                        left <= data1[678:678];
                            middle <= data2[678:678];
                            right <= data3[678:678];
                        end
                    679:
                        begin
                        left <= data1[679:679];
                            middle <= data2[679:679];
                            right <= data3[679:679];
                        end
                    680:
                        begin
                        left <= data1[680:680];
                            middle <= data2[680:680];
                            right <= data3[680:680];
                        end
                    681:
                        begin
                        left <= data1[681:681];
                            middle <= data2[681:681];
                            right <= data3[681:681];
                        end
                    682:
                        begin
                        left <= data1[682:682];
                            middle <= data2[682:682];
                            right <= data3[682:682];
                        end
                    683:
                        begin
                        left <= data1[683:683];
                            middle <= data2[683:683];
                            right <= data3[683:683];
                        end
                    684:
                        begin
                        left <= data1[684:684];
                            middle <= data2[684:684];
                            right <= data3[684:684];
                        end
                    685:
                        begin
                        left <= data1[685:685];
                            middle <= data2[685:685];
                            right <= data3[685:685];
                        end
                    686:
                        begin
                        left <= data1[686:686];
                            middle <= data2[686:686];
                            right <= data3[686:686];
                        end
                    687:
                        begin
                        left <= data1[687:687];
                            middle <= data2[687:687];
                            right <= data3[687:687];
                        end
                    688:
                        begin
                        left <= data1[688:688];
                            middle <= data2[688:688];
                            right <= data3[688:688];
                        end
                    689:
                        begin
                        left <= data1[689:689];
                            middle <= data2[689:689];
                            right <= data3[689:689];
                        end
                    690:
                        begin
                        left <= data1[690:690];
                            middle <= data2[690:690];
                            right <= data3[690:690];
                        end
                    691:
                        begin
                        left <= data1[691:691];
                            middle <= data2[691:691];
                            right <= data3[691:691];
                        end
                    692:
                        begin
                        left <= data1[692:692];
                            middle <= data2[692:692];
                            right <= data3[692:692];
                        end
                    693:
                        begin
                        left <= data1[693:693];
                            middle <= data2[693:693];
                            right <= data3[693:693];
                        end
                    694:
                        begin
                        left <= data1[694:694];
                            middle <= data2[694:694];
                            right <= data3[694:694];
                        end
                    695:
                        begin
                        left <= data1[695:695];
                            middle <= data2[695:695];
                            right <= data3[695:695];
                        end
                    696:
                        begin
                        left <= data1[696:696];
                            middle <= data2[696:696];
                            right <= data3[696:696];
                        end
                    697:
                        begin
                        left <= data1[697:697];
                            middle <= data2[697:697];
                            right <= data3[697:697];
                        end
                    698:
                        begin
                        left <= data1[698:698];
                            middle <= data2[698:698];
                            right <= data3[698:698];
                        end
                    699:
                        begin
                        left <= data1[699:699];
                            middle <= data2[699:699];
                            right <= data3[699:699];
                        end
                    700:
                        begin
                        left <= data1[700:700];
                            middle <= data2[700:700];
                            right <= data3[700:700];
                        end
                    701:
                        begin
                        left <= data1[701:701];
                            middle <= data2[701:701];
                            right <= data3[701:701];
                        end
                    702:
                        begin
                        left <= data1[702:702];
                            middle <= data2[702:702];
                            right <= data3[702:702];
                        end
                    703:
                        begin
                        left <= data1[703:703];
                            middle <= data2[703:703];
                            right <= data3[703:703];
                        end
                    704:
                        begin
                        left <= data1[704:704];
                            middle <= data2[704:704];
                            right <= data3[704:704];
                        end
                    705:
                        begin
                        left <= data1[705:705];
                            middle <= data2[705:705];
                            right <= data3[705:705];
                        end
                    706:
                        begin
                        left <= data1[706:706];
                            middle <= data2[706:706];
                            right <= data3[706:706];
                        end
                    707:
                        begin
                        left <= data1[707:707];
                            middle <= data2[707:707];
                            right <= data3[707:707];
                        end
                    708:
                        begin
                        left <= data1[708:708];
                            middle <= data2[708:708];
                            right <= data3[708:708];
                        end
                    709:
                        begin
                        left <= data1[709:709];
                            middle <= data2[709:709];
                            right <= data3[709:709];
                        end
                    710:
                        begin
                        left <= data1[710:710];
                            middle <= data2[710:710];
                            right <= data3[710:710];
                        end
                    711:
                        begin
                        left <= data1[711:711];
                            middle <= data2[711:711];
                            right <= data3[711:711];
                        end
                    712:
                        begin
                        left <= data1[712:712];
                            middle <= data2[712:712];
                            right <= data3[712:712];
                        end
                    713:
                        begin
                        left <= data1[713:713];
                            middle <= data2[713:713];
                            right <= data3[713:713];
                        end
                    714:
                        begin
                        left <= data1[714:714];
                            middle <= data2[714:714];
                            right <= data3[714:714];
                        end
                    715:
                        begin
                        left <= data1[715:715];
                            middle <= data2[715:715];
                            right <= data3[715:715];
                        end
                    716:
                        begin
                        left <= data1[716:716];
                            middle <= data2[716:716];
                            right <= data3[716:716];
                        end
                    717:
                        begin
                        left <= data1[717:717];
                            middle <= data2[717:717];
                            right <= data3[717:717];
                        end
                    718:
                        begin
                        left <= data1[718:718];
                            middle <= data2[718:718];
                            right <= data3[718:718];
                        end
                    719:
                        begin
                        left <= data1[719:719];
                            middle <= data2[719:719];
                            right <= data3[719:719];
                        end
                    720:
                        begin
                        left <= data1[720:720];
                            middle <= data2[720:720];
                            right <= data3[720:720];
                        end
                    721:
                        begin
                        left <= data1[721:721];
                            middle <= data2[721:721];
                            right <= data3[721:721];
                        end
                    722:
                        begin
                        left <= data1[722:722];
                            middle <= data2[722:722];
                            right <= data3[722:722];
                        end
                    723:
                        begin
                        left <= data1[723:723];
                            middle <= data2[723:723];
                            right <= data3[723:723];
                        end
                    724:
                        begin
                        left <= data1[724:724];
                            middle <= data2[724:724];
                            right <= data3[724:724];
                        end
                    725:
                        begin
                        left <= data1[725:725];
                            middle <= data2[725:725];
                            right <= data3[725:725];
                        end
                    726:
                        begin
                        left <= data1[726:726];
                            middle <= data2[726:726];
                            right <= data3[726:726];
                        end
                    727:
                        begin
                        left <= data1[727:727];
                            middle <= data2[727:727];
                            right <= data3[727:727];
                        end
                    728:
                        begin
                        left <= data1[728:728];
                            middle <= data2[728:728];
                            right <= data3[728:728];
                        end
                    729:
                        begin
                        left <= data1[729:729];
                            middle <= data2[729:729];
                            right <= data3[729:729];
                        end
                    730:
                        begin
                        left <= data1[730:730];
                            middle <= data2[730:730];
                            right <= data3[730:730];
                        end
                    731:
                        begin
                        left <= data1[731:731];
                            middle <= data2[731:731];
                            right <= data3[731:731];
                        end
                    732:
                        begin
                        left <= data1[732:732];
                            middle <= data2[732:732];
                            right <= data3[732:732];
                        end
                    733:
                        begin
                        left <= data1[733:733];
                            middle <= data2[733:733];
                            right <= data3[733:733];
                        end
                    734:
                        begin
                        left <= data1[734:734];
                            middle <= data2[734:734];
                            right <= data3[734:734];
                        end
                    735:
                        begin
                        left <= data1[735:735];
                            middle <= data2[735:735];
                            right <= data3[735:735];
                        end
                    736:
                        begin
                        left <= data1[736:736];
                            middle <= data2[736:736];
                            right <= data3[736:736];
                        end
                    737:
                        begin
                        left <= data1[737:737];
                            middle <= data2[737:737];
                            right <= data3[737:737];
                        end
                    738:
                        begin
                        left <= data1[738:738];
                            middle <= data2[738:738];
                            right <= data3[738:738];
                        end
                    739:
                        begin
                        left <= data1[739:739];
                            middle <= data2[739:739];
                            right <= data3[739:739];
                        end
                    740:
                        begin
                        left <= data1[740:740];
                            middle <= data2[740:740];
                            right <= data3[740:740];
                        end
                    741:
                        begin
                        left <= data1[741:741];
                            middle <= data2[741:741];
                            right <= data3[741:741];
                        end
                    742:
                        begin
                        left <= data1[742:742];
                            middle <= data2[742:742];
                            right <= data3[742:742];
                        end
                    743:
                        begin
                        left <= data1[743:743];
                            middle <= data2[743:743];
                            right <= data3[743:743];
                        end
                    744:
                        begin
                        left <= data1[744:744];
                            middle <= data2[744:744];
                            right <= data3[744:744];
                        end
                    745:
                        begin
                        left <= data1[745:745];
                            middle <= data2[745:745];
                            right <= data3[745:745];
                        end
                    746:
                        begin
                        left <= data1[746:746];
                            middle <= data2[746:746];
                            right <= data3[746:746];
                        end
                    747:
                        begin
                        left <= data1[747:747];
                            middle <= data2[747:747];
                            right <= data3[747:747];
                        end
                    748:
                        begin
                        left <= data1[748:748];
                            middle <= data2[748:748];
                            right <= data3[748:748];
                        end
                    749:
                        begin
                        left <= data1[749:749];
                            middle <= data2[749:749];
                            right <= data3[749:749];
                        end
                    750:
                        begin
                        left <= data1[750:750];
                            middle <= data2[750:750];
                            right <= data3[750:750];
                        end
                    751:
                        begin
                        left <= data1[751:751];
                            middle <= data2[751:751];
                            right <= data3[751:751];
                        end
                    752:
                        begin
                        left <= data1[752:752];
                            middle <= data2[752:752];
                            right <= data3[752:752];
                        end
                    753:
                        begin
                        left <= data1[753:753];
                            middle <= data2[753:753];
                            right <= data3[753:753];
                        end
                    754:
                        begin
                        left <= data1[754:754];
                            middle <= data2[754:754];
                            right <= data3[754:754];
                        end
                    755:
                        begin
                        left <= data1[755:755];
                            middle <= data2[755:755];
                            right <= data3[755:755];
                        end
                    756:
                        begin
                        left <= data1[756:756];
                            middle <= data2[756:756];
                            right <= data3[756:756];
                        end
                    757:
                        begin
                        left <= data1[757:757];
                            middle <= data2[757:757];
                            right <= data3[757:757];
                        end
                    758:
                        begin
                        left <= data1[758:758];
                            middle <= data2[758:758];
                            right <= data3[758:758];
                        end
                    759:
                        begin
                        left <= data1[759:759];
                            middle <= data2[759:759];
                            right <= data3[759:759];
                        end
                    760:
                        begin
                        left <= data1[760:760];
                            middle <= data2[760:760];
                            right <= data3[760:760];
                        end
                    761:
                        begin
                        left <= data1[761:761];
                            middle <= data2[761:761];
                            right <= data3[761:761];
                        end
                    762:
                        begin
                        left <= data1[762:762];
                            middle <= data2[762:762];
                            right <= data3[762:762];
                        end
                    763:
                        begin
                        left <= data1[763:763];
                            middle <= data2[763:763];
                            right <= data3[763:763];
                        end
                    764:
                        begin
                        left <= data1[764:764];
                            middle <= data2[764:764];
                            right <= data3[764:764];
                        end
                    765:
                        begin
                        left <= data1[765:765];
                            middle <= data2[765:765];
                            right <= data3[765:765];
                        end
                    766:
                        begin
                        left <= data1[766:766];
                            middle <= data2[766:766];
                            right <= data3[766:766];
                        end
                    767:
                        begin
                        left <= data1[767:767];
                            middle <= data2[767:767];
                            right <= data3[767:767];
                        end
                    768:
                        begin
                        left <= data1[768:768];
                            middle <= data2[768:768];
                            right <= data3[768:768];
                        end
                    769:
                        begin
                        left <= data1[769:769];
                            middle <= data2[769:769];
                            right <= data3[769:769];
                        end
                    770:
                        begin
                        left <= data1[770:770];
                            middle <= data2[770:770];
                            right <= data3[770:770];
                        end
                    771:
                        begin
                        left <= data1[771:771];
                            middle <= data2[771:771];
                            right <= data3[771:771];
                        end
                    772:
                        begin
                        left <= data1[772:772];
                            middle <= data2[772:772];
                            right <= data3[772:772];
                        end
                    773:
                        begin
                        left <= data1[773:773];
                            middle <= data2[773:773];
                            right <= data3[773:773];
                        end
                    774:
                        begin
                        left <= data1[774:774];
                            middle <= data2[774:774];
                            right <= data3[774:774];
                        end
                    775:
                        begin
                        left <= data1[775:775];
                            middle <= data2[775:775];
                            right <= data3[775:775];
                        end
                    776:
                        begin
                        left <= data1[776:776];
                            middle <= data2[776:776];
                            right <= data3[776:776];
                        end
                    777:
                        begin
                        left <= data1[777:777];
                            middle <= data2[777:777];
                            right <= data3[777:777];
                        end
                    778:
                        begin
                        left <= data1[778:778];
                            middle <= data2[778:778];
                            right <= data3[778:778];
                        end
                    779:
                        begin
                        left <= data1[779:779];
                            middle <= data2[779:779];
                            right <= data3[779:779];
                        end
                    780:
                        begin
                        left <= data1[780:780];
                            middle <= data2[780:780];
                            right <= data3[780:780];
                        end
                    781:
                        begin
                        left <= data1[781:781];
                            middle <= data2[781:781];
                            right <= data3[781:781];
                        end
                    782:
                        begin
                        left <= data1[782:782];
                            middle <= data2[782:782];
                            right <= data3[782:782];
                        end
                    783:
                        begin
                        left <= data1[783:783];
                            middle <= data2[783:783];
                            right <= data3[783:783];
                        end
                    784:
                        begin
                        left <= data1[784:784];
                            middle <= data2[784:784];
                            right <= data3[784:784];
                        end
                    785:
                        begin
                        left <= data1[785:785];
                            middle <= data2[785:785];
                            right <= data3[785:785];
                        end
                    786:
                        begin
                        left <= data1[786:786];
                            middle <= data2[786:786];
                            right <= data3[786:786];
                        end
                    787:
                        begin
                        left <= data1[787:787];
                            middle <= data2[787:787];
                            right <= data3[787:787];
                        end
                    788:
                        begin
                        left <= data1[788:788];
                            middle <= data2[788:788];
                            right <= data3[788:788];
                        end
                    789:
                        begin
                        left <= data1[789:789];
                            middle <= data2[789:789];
                            right <= data3[789:789];
                        end
                    790:
                        begin
                        left <= data1[790:790];
                            middle <= data2[790:790];
                            right <= data3[790:790];
                        end
                    791:
                        begin
                        left <= data1[791:791];
                            middle <= data2[791:791];
                            right <= data3[791:791];
                        end
                    792:
                        begin
                        left <= data1[792:792];
                            middle <= data2[792:792];
                            right <= data3[792:792];
                        end
                    793:
                        begin
                        left <= data1[793:793];
                            middle <= data2[793:793];
                            right <= data3[793:793];
                        end
                    794:
                        begin
                        left <= data1[794:794];
                            middle <= data2[794:794];
                            right <= data3[794:794];
                        end
                    795:
                        begin
                        left <= data1[795:795];
                            middle <= data2[795:795];
                            right <= data3[795:795];
                        end
                    796:
                        begin
                        left <= data1[796:796];
                            middle <= data2[796:796];
                            right <= data3[796:796];
                        end
                    797:
                        begin
                        left <= data1[797:797];
                            middle <= data2[797:797];
                            right <= data3[797:797];
                        end
                    798:
                        begin
                        left <= data1[798:798];
                            middle <= data2[798:798];
                            right <= data3[798:798];
                        end
                    799:
                        begin
                        left <= data1[799:799];
                            middle <= data2[799:799];
                            right <= data3[799:799];
                        end
                    800:
                        begin
                        left <= data1[800:800];
                            middle <= data2[800:800];
                            right <= data3[800:800];
                        end
                    801:
                        begin
                        left <= data1[801:801];
                            middle <= data2[801:801];
                            right <= data3[801:801];
                        end
                    802:
                        begin
                        left <= data1[802:802];
                            middle <= data2[802:802];
                            right <= data3[802:802];
                        end
                    803:
                        begin
                        left <= data1[803:803];
                            middle <= data2[803:803];
                            right <= data3[803:803];
                        end
                    804:
                        begin
                        left <= data1[804:804];
                            middle <= data2[804:804];
                            right <= data3[804:804];
                        end
                    805:
                        begin
                        left <= data1[805:805];
                            middle <= data2[805:805];
                            right <= data3[805:805];
                        end
                    806:
                        begin
                        left <= data1[806:806];
                            middle <= data2[806:806];
                            right <= data3[806:806];
                        end
                    807:
                        begin
                        left <= data1[807:807];
                            middle <= data2[807:807];
                            right <= data3[807:807];
                        end
                    808:
                        begin
                        left <= data1[808:808];
                            middle <= data2[808:808];
                            right <= data3[808:808];
                        end
                    809:
                        begin
                        left <= data1[809:809];
                            middle <= data2[809:809];
                            right <= data3[809:809];
                        end
                    810:
                        begin
                        left <= data1[810:810];
                            middle <= data2[810:810];
                            right <= data3[810:810];
                        end
                    811:
                        begin
                        left <= data1[811:811];
                            middle <= data2[811:811];
                            right <= data3[811:811];
                        end
                    812:
                        begin
                        left <= data1[812:812];
                            middle <= data2[812:812];
                            right <= data3[812:812];
                        end
                    813:
                        begin
                        left <= data1[813:813];
                            middle <= data2[813:813];
                            right <= data3[813:813];
                        end
                    814:
                        begin
                        left <= data1[814:814];
                            middle <= data2[814:814];
                            right <= data3[814:814];
                        end
                    815:
                        begin
                        left <= data1[815:815];
                            middle <= data2[815:815];
                            right <= data3[815:815];
                        end
                    816:
                        begin
                        left <= data1[816:816];
                            middle <= data2[816:816];
                            right <= data3[816:816];
                        end
                    817:
                        begin
                        left <= data1[817:817];
                            middle <= data2[817:817];
                            right <= data3[817:817];
                        end
                    818:
                        begin
                        left <= data1[818:818];
                            middle <= data2[818:818];
                            right <= data3[818:818];
                        end
                    819:
                        begin
                        left <= data1[819:819];
                            middle <= data2[819:819];
                            right <= data3[819:819];
                        end
                    820:
                        begin
                        left <= data1[820:820];
                            middle <= data2[820:820];
                            right <= data3[820:820];
                        end
                    821:
                        begin
                        left <= data1[821:821];
                            middle <= data2[821:821];
                            right <= data3[821:821];
                        end
                    822:
                        begin
                        left <= data1[822:822];
                            middle <= data2[822:822];
                            right <= data3[822:822];
                        end
                    823:
                        begin
                        left <= data1[823:823];
                            middle <= data2[823:823];
                            right <= data3[823:823];
                        end
                    824:
                        begin
                        left <= data1[824:824];
                            middle <= data2[824:824];
                            right <= data3[824:824];
                        end
                    825:
                        begin
                        left <= data1[825:825];
                            middle <= data2[825:825];
                            right <= data3[825:825];
                        end
                    826:
                        begin
                        left <= data1[826:826];
                            middle <= data2[826:826];
                            right <= data3[826:826];
                        end
                    827:
                        begin
                        left <= data1[827:827];
                            middle <= data2[827:827];
                            right <= data3[827:827];
                        end
                    828:
                        begin
                        left <= data1[828:828];
                            middle <= data2[828:828];
                            right <= data3[828:828];
                        end
                    829:
                        begin
                        left <= data1[829:829];
                            middle <= data2[829:829];
                            right <= data3[829:829];
                        end
                    830:
                        begin
                        left <= data1[830:830];
                            middle <= data2[830:830];
                            right <= data3[830:830];
                        end
                    831:
                        begin
                        left <= data1[831:831];
                            middle <= data2[831:831];
                            right <= data3[831:831];
                        end
                    832:
                        begin
                        left <= data1[832:832];
                            middle <= data2[832:832];
                            right <= data3[832:832];
                        end
                    833:
                        begin
                        left <= data1[833:833];
                            middle <= data2[833:833];
                            right <= data3[833:833];
                        end
                    834:
                        begin
                        left <= data1[834:834];
                            middle <= data2[834:834];
                            right <= data3[834:834];
                        end
                    835:
                        begin
                        left <= data1[835:835];
                            middle <= data2[835:835];
                            right <= data3[835:835];
                        end
                    836:
                        begin
                        left <= data1[836:836];
                            middle <= data2[836:836];
                            right <= data3[836:836];
                        end
                    837:
                        begin
                        left <= data1[837:837];
                            middle <= data2[837:837];
                            right <= data3[837:837];
                        end
                    838:
                        begin
                        left <= data1[838:838];
                            middle <= data2[838:838];
                            right <= data3[838:838];
                        end
                    839:
                        begin
                        left <= data1[839:839];
                            middle <= data2[839:839];
                            right <= data3[839:839];
                        end
                    840:
                        begin
                        left <= data1[840:840];
                            middle <= data2[840:840];
                            right <= data3[840:840];
                        end
                    841:
                        begin
                        left <= data1[841:841];
                            middle <= data2[841:841];
                            right <= data3[841:841];
                        end
                    842:
                        begin
                        left <= data1[842:842];
                            middle <= data2[842:842];
                            right <= data3[842:842];
                        end
                    843:
                        begin
                        left <= data1[843:843];
                            middle <= data2[843:843];
                            right <= data3[843:843];
                        end
                    844:
                        begin
                        left <= data1[844:844];
                            middle <= data2[844:844];
                            right <= data3[844:844];
                        end
                    845:
                        begin
                        left <= data1[845:845];
                            middle <= data2[845:845];
                            right <= data3[845:845];
                        end
                    846:
                        begin
                        left <= data1[846:846];
                            middle <= data2[846:846];
                            right <= data3[846:846];
                        end
                    847:
                        begin
                        left <= data1[847:847];
                            middle <= data2[847:847];
                            right <= data3[847:847];
                        end
                    848:
                        begin
                        left <= data1[848:848];
                            middle <= data2[848:848];
                            right <= data3[848:848];
                        end
                    849:
                        begin
                        left <= data1[849:849];
                            middle <= data2[849:849];
                            right <= data3[849:849];
                        end
                    850:
                        begin
                        left <= data1[850:850];
                            middle <= data2[850:850];
                            right <= data3[850:850];
                        end
                    851:
                        begin
                        left <= data1[851:851];
                            middle <= data2[851:851];
                            right <= data3[851:851];
                        end
                    852:
                        begin
                        left <= data1[852:852];
                            middle <= data2[852:852];
                            right <= data3[852:852];
                        end
                    853:
                        begin
                        left <= data1[853:853];
                            middle <= data2[853:853];
                            right <= data3[853:853];
                        end
                    854:
                        begin
                        left <= data1[854:854];
                            middle <= data2[854:854];
                            right <= data3[854:854];
                        end
                    855:
                        begin
                        left <= data1[855:855];
                            middle <= data2[855:855];
                            right <= data3[855:855];
                        end
                    856:
                        begin
                        left <= data1[856:856];
                            middle <= data2[856:856];
                            right <= data3[856:856];
                        end
                    857:
                        begin
                        left <= data1[857:857];
                            middle <= data2[857:857];
                            right <= data3[857:857];
                        end
                    858:
                        begin
                        left <= data1[858:858];
                            middle <= data2[858:858];
                            right <= data3[858:858];
                        end
                    859:
                        begin
                        left <= data1[859:859];
                            middle <= data2[859:859];
                            right <= data3[859:859];
                        end
                    860:
                        begin
                        left <= data1[860:860];
                            middle <= data2[860:860];
                            right <= data3[860:860];
                        end
                    861:
                        begin
                        left <= data1[861:861];
                            middle <= data2[861:861];
                            right <= data3[861:861];
                        end
                    862:
                        begin
                        left <= data1[862:862];
                            middle <= data2[862:862];
                            right <= data3[862:862];
                        end
                    863:
                        begin
                        left <= data1[863:863];
                            middle <= data2[863:863];
                            right <= data3[863:863];
                        end
                    864:
                        begin
                        left <= data1[864:864];
                            middle <= data2[864:864];
                            right <= data3[864:864];
                        end
                    865:
                        begin
                        left <= data1[865:865];
                            middle <= data2[865:865];
                            right <= data3[865:865];
                        end
                    866:
                        begin
                        left <= data1[866:866];
                            middle <= data2[866:866];
                            right <= data3[866:866];
                        end
                    867:
                        begin
                        left <= data1[867:867];
                            middle <= data2[867:867];
                            right <= data3[867:867];
                        end
                    868:
                        begin
                        left <= data1[868:868];
                            middle <= data2[868:868];
                            right <= data3[868:868];
                        end
                    869:
                        begin
                        left <= data1[869:869];
                            middle <= data2[869:869];
                            right <= data3[869:869];
                        end
                    870:
                        begin
                        left <= data1[870:870];
                            middle <= data2[870:870];
                            right <= data3[870:870];
                        end
                    871:
                        begin
                        left <= data1[871:871];
                            middle <= data2[871:871];
                            right <= data3[871:871];
                        end
                    872:
                        begin
                        left <= data1[872:872];
                            middle <= data2[872:872];
                            right <= data3[872:872];
                        end
                    873:
                        begin
                        left <= data1[873:873];
                            middle <= data2[873:873];
                            right <= data3[873:873];
                        end
                    874:
                        begin
                        left <= data1[874:874];
                            middle <= data2[874:874];
                            right <= data3[874:874];
                        end
                    875:
                        begin
                        left <= data1[875:875];
                            middle <= data2[875:875];
                            right <= data3[875:875];
                        end
                    876:
                        begin
                        left <= data1[876:876];
                            middle <= data2[876:876];
                            right <= data3[876:876];
                        end
                    877:
                        begin
                        left <= data1[877:877];
                            middle <= data2[877:877];
                            right <= data3[877:877];
                        end
                    878:
                        begin
                        left <= data1[878:878];
                            middle <= data2[878:878];
                            right <= data3[878:878];
                        end
                    879:
                        begin
                        left <= data1[879:879];
                            middle <= data2[879:879];
                            right <= data3[879:879];
                        end
                    880:
                        begin
                        left <= data1[880:880];
                            middle <= data2[880:880];
                            right <= data3[880:880];
                        end
                    881:
                        begin
                        left <= data1[881:881];
                            middle <= data2[881:881];
                            right <= data3[881:881];
                        end
                    882:
                        begin
                        left <= data1[882:882];
                            middle <= data2[882:882];
                            right <= data3[882:882];
                        end
                    883:
                        begin
                        left <= data1[883:883];
                            middle <= data2[883:883];
                            right <= data3[883:883];
                        end
                    884:
                        begin
                        left <= data1[884:884];
                            middle <= data2[884:884];
                            right <= data3[884:884];
                        end
                    885:
                        begin
                        left <= data1[885:885];
                            middle <= data2[885:885];
                            right <= data3[885:885];
                        end
                    886:
                        begin
                        left <= data1[886:886];
                            middle <= data2[886:886];
                            right <= data3[886:886];
                        end
                    887:
                        begin
                        left <= data1[887:887];
                            middle <= data2[887:887];
                            right <= data3[887:887];
                        end
                    888:
                        begin
                        left <= data1[888:888];
                            middle <= data2[888:888];
                            right <= data3[888:888];
                        end
                    889:
                        begin
                        left <= data1[889:889];
                            middle <= data2[889:889];
                            right <= data3[889:889];
                        end
                    890:
                        begin
                        left <= data1[890:890];
                            middle <= data2[890:890];
                            right <= data3[890:890];
                        end
                    891:
                        begin
                        left <= data1[891:891];
                            middle <= data2[891:891];
                            right <= data3[891:891];
                        end
                    892:
                        begin
                        left <= data1[892:892];
                            middle <= data2[892:892];
                            right <= data3[892:892];
                        end
                    893:
                        begin
                        left <= data1[893:893];
                            middle <= data2[893:893];
                            right <= data3[893:893];
                        end
                    894:
                        begin
                        left <= data1[894:894];
                            middle <= data2[894:894];
                            right <= data3[894:894];
                        end
                    895:
                        begin
                        left <= data1[895:895];
                            middle <= data2[895:895];
                            right <= data3[895:895];
                        end
                    896:
                        begin
                        left <= data1[896:896];
                            middle <= data2[896:896];
                            right <= data3[896:896];
                        end
                    897:
                        begin
                        left <= data1[897:897];
                            middle <= data2[897:897];
                            right <= data3[897:897];
                        end
                    898:
                        begin
                        left <= data1[898:898];
                            middle <= data2[898:898];
                            right <= data3[898:898];
                        end
                    899:
                        begin
                        left <= data1[899:899];
                            middle <= data2[899:899];
                            right <= data3[899:899];
                        end
                    900:
                        begin
                        left <= data1[900:900];
                            middle <= data2[900:900];
                            right <= data3[900:900];
                        end
                    901:
                        begin
                        left <= data1[901:901];
                            middle <= data2[901:901];
                            right <= data3[901:901];
                        end
                    902:
                        begin
                        left <= data1[902:902];
                            middle <= data2[902:902];
                            right <= data3[902:902];
                        end
                    903:
                        begin
                        left <= data1[903:903];
                            middle <= data2[903:903];
                            right <= data3[903:903];
                        end
                    904:
                        begin
                        left <= data1[904:904];
                            middle <= data2[904:904];
                            right <= data3[904:904];
                        end
                    905:
                        begin
                        left <= data1[905:905];
                            middle <= data2[905:905];
                            right <= data3[905:905];
                        end
                    906:
                        begin
                        left <= data1[906:906];
                            middle <= data2[906:906];
                            right <= data3[906:906];
                        end
                    907:
                        begin
                        left <= data1[907:907];
                            middle <= data2[907:907];
                            right <= data3[907:907];
                        end
                    908:
                        begin
                        left <= data1[908:908];
                            middle <= data2[908:908];
                            right <= data3[908:908];
                        end
                    909:
                        begin
                        left <= data1[909:909];
                            middle <= data2[909:909];
                            right <= data3[909:909];
                        end
                    910:
                        begin
                        left <= data1[910:910];
                            middle <= data2[910:910];
                            right <= data3[910:910];
                        end
                    911:
                        begin
                        left <= data1[911:911];
                            middle <= data2[911:911];
                            right <= data3[911:911];
                        end
                    912:
                        begin
                        left <= data1[912:912];
                            middle <= data2[912:912];
                            right <= data3[912:912];
                        end
                    913:
                        begin
                        left <= data1[913:913];
                            middle <= data2[913:913];
                            right <= data3[913:913];
                        end
                    914:
                        begin
                        left <= data1[914:914];
                            middle <= data2[914:914];
                            right <= data3[914:914];
                        end
                    915:
                        begin
                        left <= data1[915:915];
                            middle <= data2[915:915];
                            right <= data3[915:915];
                        end
                    916:
                        begin
                        left <= data1[916:916];
                            middle <= data2[916:916];
                            right <= data3[916:916];
                        end
                    917:
                        begin
                        left <= data1[917:917];
                            middle <= data2[917:917];
                            right <= data3[917:917];
                        end
                    918:
                        begin
                        left <= data1[918:918];
                            middle <= data2[918:918];
                            right <= data3[918:918];
                        end
                    919:
                        begin
                        left <= data1[919:919];
                            middle <= data2[919:919];
                            right <= data3[919:919];
                        end
                    920:
                        begin
                        left <= data1[920:920];
                            middle <= data2[920:920];
                            right <= data3[920:920];
                        end
                    921:
                        begin
                        left <= data1[921:921];
                            middle <= data2[921:921];
                            right <= data3[921:921];
                        end
                    922:
                        begin
                        left <= data1[922:922];
                            middle <= data2[922:922];
                            right <= data3[922:922];
                        end
                    923:
                        begin
                        left <= data1[923:923];
                            middle <= data2[923:923];
                            right <= data3[923:923];
                        end
                    924:
                        begin
                        left <= data1[924:924];
                            middle <= data2[924:924];
                            right <= data3[924:924];
                        end
                    925:
                        begin
                        left <= data1[925:925];
                            middle <= data2[925:925];
                            right <= data3[925:925];
                        end
                    926:
                        begin
                        left <= data1[926:926];
                            middle <= data2[926:926];
                            right <= data3[926:926];
                        end
                    927:
                        begin
                        left <= data1[927:927];
                            middle <= data2[927:927];
                            right <= data3[927:927];
                        end
                    928:
                        begin
                        left <= data1[928:928];
                            middle <= data2[928:928];
                            right <= data3[928:928];
                        end
                    929:
                        begin
                        left <= data1[929:929];
                            middle <= data2[929:929];
                            right <= data3[929:929];
                        end
                    930:
                        begin
                        left <= data1[930:930];
                            middle <= data2[930:930];
                            right <= data3[930:930];
                        end
                    931:
                        begin
                        left <= data1[931:931];
                            middle <= data2[931:931];
                            right <= data3[931:931];
                        end
                    932:
                        begin
                        left <= data1[932:932];
                            middle <= data2[932:932];
                            right <= data3[932:932];
                        end
                    933:
                        begin
                        left <= data1[933:933];
                            middle <= data2[933:933];
                            right <= data3[933:933];
                        end
                    934:
                        begin
                        left <= data1[934:934];
                            middle <= data2[934:934];
                            right <= data3[934:934];
                        end
                    935:
                        begin
                        left <= data1[935:935];
                            middle <= data2[935:935];
                            right <= data3[935:935];
                        end
                    936:
                        begin
                        left <= data1[936:936];
                            middle <= data2[936:936];
                            right <= data3[936:936];
                        end
                    937:
                        begin
                        left <= data1[937:937];
                            middle <= data2[937:937];
                            right <= data3[937:937];
                        end
                    938:
                        begin
                        left <= data1[938:938];
                            middle <= data2[938:938];
                            right <= data3[938:938];
                        end
                    939:
                        begin
                        left <= data1[939:939];
                            middle <= data2[939:939];
                            right <= data3[939:939];
                        end
                    940:
                        begin
                        left <= data1[940:940];
                            middle <= data2[940:940];
                            right <= data3[940:940];
                        end
                    941:
                        begin
                        left <= data1[941:941];
                            middle <= data2[941:941];
                            right <= data3[941:941];
                        end
                    942:
                        begin
                        left <= data1[942:942];
                            middle <= data2[942:942];
                            right <= data3[942:942];
                        end
                    943:
                        begin
                        left <= data1[943:943];
                            middle <= data2[943:943];
                            right <= data3[943:943];
                        end
                    944:
                        begin
                        left <= data1[944:944];
                            middle <= data2[944:944];
                            right <= data3[944:944];
                        end
                    945:
                        begin
                        left <= data1[945:945];
                            middle <= data2[945:945];
                            right <= data3[945:945];
                        end
                    946:
                        begin
                        left <= data1[946:946];
                            middle <= data2[946:946];
                            right <= data3[946:946];
                        end
                    947:
                        begin
                        left <= data1[947:947];
                            middle <= data2[947:947];
                            right <= data3[947:947];
                        end
                    948:
                        begin
                        left <= data1[948:948];
                            middle <= data2[948:948];
                            right <= data3[948:948];
                        end
                    949:
                        begin
                        left <= data1[949:949];
                            middle <= data2[949:949];
                            right <= data3[949:949];
                        end
                    950:
                        begin
                        left <= data1[950:950];
                            middle <= data2[950:950];
                            right <= data3[950:950];
                        end
                    951:
                        begin
                        left <= data1[951:951];
                            middle <= data2[951:951];
                            right <= data3[951:951];
                        end
                    952:
                        begin
                        left <= data1[952:952];
                            middle <= data2[952:952];
                            right <= data3[952:952];
                        end
                    953:
                        begin
                        left <= data1[953:953];
                            middle <= data2[953:953];
                            right <= data3[953:953];
                        end
                    954:
                        begin
                        left <= data1[954:954];
                            middle <= data2[954:954];
                            right <= data3[954:954];
                        end
                    955:
                        begin
                        left <= data1[955:955];
                            middle <= data2[955:955];
                            right <= data3[955:955];
                        end
                    956:
                        begin
                        left <= data1[956:956];
                            middle <= data2[956:956];
                            right <= data3[956:956];
                        end
                    957:
                        begin
                        left <= data1[957:957];
                            middle <= data2[957:957];
                            right <= data3[957:957];
                        end
                    958:
                        begin
                        left <= data1[958:958];
                            middle <= data2[958:958];
                            right <= data3[958:958];
                        end
                    959:
                        begin
                        left <= data1[959:959];
                            middle <= data2[959:959];
                            right <= data3[959:959];
                        end
                    960:
                        begin
                        left <= data1[960:960];
                            middle <= data2[960:960];
                            right <= data3[960:960];
                        end
                    961:
                        begin
                        left <= data1[961:961];
                            middle <= data2[961:961];
                            right <= data3[961:961];
                        end
                    962:
                        begin
                        left <= data1[962:962];
                            middle <= data2[962:962];
                            right <= data3[962:962];
                        end
                    963:
                        begin
                        left <= data1[963:963];
                            middle <= data2[963:963];
                            right <= data3[963:963];
                        end
                    964:
                        begin
                        left <= data1[964:964];
                            middle <= data2[964:964];
                            right <= data3[964:964];
                        end
                    965:
                        begin
                        left <= data1[965:965];
                            middle <= data2[965:965];
                            right <= data3[965:965];
                        end
                    966:
                        begin
                        left <= data1[966:966];
                            middle <= data2[966:966];
                            right <= data3[966:966];
                        end
                    967:
                        begin
                        left <= data1[967:967];
                            middle <= data2[967:967];
                            right <= data3[967:967];
                        end
                    968:
                        begin
                        left <= data1[968:968];
                            middle <= data2[968:968];
                            right <= data3[968:968];
                        end
                    969:
                        begin
                        left <= data1[969:969];
                            middle <= data2[969:969];
                            right <= data3[969:969];
                        end
                    970:
                        begin
                        left <= data1[970:970];
                            middle <= data2[970:970];
                            right <= data3[970:970];
                        end
                    971:
                        begin
                        left <= data1[971:971];
                            middle <= data2[971:971];
                            right <= data3[971:971];
                        end
                    972:
                        begin
                        left <= data1[972:972];
                            middle <= data2[972:972];
                            right <= data3[972:972];
                        end
                    973:
                        begin
                        left <= data1[973:973];
                            middle <= data2[973:973];
                            right <= data3[973:973];
                        end
                    974:
                        begin
                        left <= data1[974:974];
                            middle <= data2[974:974];
                            right <= data3[974:974];
                        end
                    975:
                        begin
                        left <= data1[975:975];
                            middle <= data2[975:975];
                            right <= data3[975:975];
                        end
                    976:
                        begin
                        left <= data1[976:976];
                            middle <= data2[976:976];
                            right <= data3[976:976];
                        end
                    977:
                        begin
                        left <= data1[977:977];
                            middle <= data2[977:977];
                            right <= data3[977:977];
                        end
                    978:
                        begin
                        left <= data1[978:978];
                            middle <= data2[978:978];
                            right <= data3[978:978];
                        end
                    979:
                        begin
                        left <= data1[979:979];
                            middle <= data2[979:979];
                            right <= data3[979:979];
                        end
                    980:
                        begin
                        left <= data1[980:980];
                            middle <= data2[980:980];
                            right <= data3[980:980];
                        end
                    981:
                        begin
                        left <= data1[981:981];
                            middle <= data2[981:981];
                            right <= data3[981:981];
                        end
                    982:
                        begin
                        left <= data1[982:982];
                            middle <= data2[982:982];
                            right <= data3[982:982];
                        end
                    983:
                        begin
                        left <= data1[983:983];
                            middle <= data2[983:983];
                            right <= data3[983:983];
                        end
                    984:
                        begin
                        left <= data1[984:984];
                            middle <= data2[984:984];
                            right <= data3[984:984];
                        end
                    985:
                        begin
                        left <= data1[985:985];
                            middle <= data2[985:985];
                            right <= data3[985:985];
                        end
                    986:
                        begin
                        left <= data1[986:986];
                            middle <= data2[986:986];
                            right <= data3[986:986];
                        end
                    987:
                        begin
                        left <= data1[987:987];
                            middle <= data2[987:987];
                            right <= data3[987:987];
                        end
                    988:
                        begin
                        left <= data1[988:988];
                            middle <= data2[988:988];
                            right <= data3[988:988];
                        end
                    989:
                        begin
                        left <= data1[989:989];
                            middle <= data2[989:989];
                            right <= data3[989:989];
                        end
                    990:
                        begin
                        left <= data1[990:990];
                            middle <= data2[990:990];
                            right <= data3[990:990];
                        end
                    991:
                        begin
                        left <= data1[991:991];
                            middle <= data2[991:991];
                            right <= data3[991:991];
                        end
                    992:
                        begin
                        left <= data1[992:992];
                            middle <= data2[992:992];
                            right <= data3[992:992];
                        end
                    993:
                        begin
                        left <= data1[993:993];
                            middle <= data2[993:993];
                            right <= data3[993:993];
                        end
                    994:
                        begin
                        left <= data1[994:994];
                            middle <= data2[994:994];
                            right <= data3[994:994];
                        end
                    995:
                        begin
                        left <= data1[995:995];
                            middle <= data2[995:995];
                            right <= data3[995:995];
                        end
                    996:
                        begin
                        left <= data1[996:996];
                            middle <= data2[996:996];
                            right <= data3[996:996];
                        end
                    997:
                        begin
                        left <= data1[997:997];
                            middle <= data2[997:997];
                            right <= data3[997:997];
                        end
                    998:
                        begin
                        left <= data1[998:998];
                            middle <= data2[998:998];
                            right <= data3[998:998];
                        end
                    999:
                        begin
                        left <= data1[999:999];
                            middle <= data2[999:999];
                            right <= data3[999:999];
                        end
                    1000:
                        begin
                        left <= data1[1000:1000];
                            middle <= data2[1000:1000];
                            right <= data3[1000:1000];
                        end
                    1001:
                        begin
                        left <= data1[1001:1001];
                            middle <= data2[1001:1001];
                            right <= data3[1001:1001];
                        end
                    1002:
                        begin
                        left <= data1[1002:1002];
                            middle <= data2[1002:1002];
                            right <= data3[1002:1002];
                        end
                    1003:
                        begin
                        left <= data1[1003:1003];
                            middle <= data2[1003:1003];
                            right <= data3[1003:1003];
                        end
                    1004:
                        begin
                        left <= data1[1004:1004];
                            middle <= data2[1004:1004];
                            right <= data3[1004:1004];
                        end
                    1005:
                        begin
                        left <= data1[1005:1005];
                            middle <= data2[1005:1005];
                            right <= data3[1005:1005];
                        end
                    1006:
                        begin
                        left <= data1[1006:1006];
                            middle <= data2[1006:1006];
                            right <= data3[1006:1006];
                        end
                    1007:
                        begin
                        left <= data1[1007:1007];
                            middle <= data2[1007:1007];
                            right <= data3[1007:1007];
                        end
                    1008:
                        begin
                        left <= data1[1008:1008];
                            middle <= data2[1008:1008];
                            right <= data3[1008:1008];
                        end
                    1009:
                        begin
                        left <= data1[1009:1009];
                            middle <= data2[1009:1009];
                            right <= data3[1009:1009];
                        end
                    1010:
                        begin
                        left <= data1[1010:1010];
                            middle <= data2[1010:1010];
                            right <= data3[1010:1010];
                        end
                    1011:
                        begin
                        left <= data1[1011:1011];
                            middle <= data2[1011:1011];
                            right <= data3[1011:1011];
                        end
                    1012:
                        begin
                        left <= data1[1012:1012];
                            middle <= data2[1012:1012];
                            right <= data3[1012:1012];
                        end
                    1013:
                        begin
                        left <= data1[1013:1013];
                            middle <= data2[1013:1013];
                            right <= data3[1013:1013];
                        end
                    1014:
                        begin
                        left <= data1[1014:1014];
                            middle <= data2[1014:1014];
                            right <= data3[1014:1014];
                        end
                    1015:
                        begin
                        left <= data1[1015:1015];
                            middle <= data2[1015:1015];
                            right <= data3[1015:1015];
                        end
                    1016:
                        begin
                        left <= data1[1016:1016];
                            middle <= data2[1016:1016];
                            right <= data3[1016:1016];
                        end
                    1017:
                        begin
                        left <= data1[1017:1017];
                            middle <= data2[1017:1017];
                            right <= data3[1017:1017];
                        end
                    1018:
                        begin
                        left <= data1[1018:1018];
                            middle <= data2[1018:1018];
                            right <= data3[1018:1018];
                        end
                    1019:
                        begin
                        left <= data1[1019:1019];
                            middle <= data2[1019:1019];
                            right <= data3[1019:1019];
                        end
                    1020:
                        begin
                        left <= data1[1020:1020];
                            middle <= data2[1020:1020];
                            right <= data3[1020:1020];
                        end
                    1021:
                        begin
                        left <= data1[1021:1021];
                            middle <= data2[1021:1021];
                            right <= data3[1021:1021];
                        end
                    1022:
                        begin
                        left <= data1[1022:1022];
                            middle <= data2[1022:1022];
                            right <= data3[1022:1022];
                        end
                    1023:
                        begin
                        left <= data1[1023:1023];
                            middle <= data2[1023:1023];
                            right <= data3[1023:1023];
                        end
                    1024:
                        begin
                        left <= data1[1024:1024];
                            middle <= data2[1024:1024];
                            right <= data3[1024:1024];
                        end
                    1025:
                        begin
                        left <= data1[1025:1025];
                            middle <= data2[1025:1025];
                            right <= data3[1025:1025];
                        end
                    1026:
                        begin
                        left <= data1[1026:1026];
                            middle <= data2[1026:1026];
                            right <= data3[1026:1026];
                        end
                    1027:
                        begin
                        left <= data1[1027:1027];
                            middle <= data2[1027:1027];
                            right <= data3[1027:1027];
                        end
                    1028:
                        begin
                        left <= data1[1028:1028];
                            middle <= data2[1028:1028];
                            right <= data3[1028:1028];
                        end
                    1029:
                        begin
                        left <= data1[1029:1029];
                            middle <= data2[1029:1029];
                            right <= data3[1029:1029];
                        end
                    1030:
                        begin
                        left <= data1[1030:1030];
                            middle <= data2[1030:1030];
                            right <= data3[1030:1030];
                        end
                    1031:
                        begin
                        left <= data1[1031:1031];
                            middle <= data2[1031:1031];
                            right <= data3[1031:1031];
                        end
                    1032:
                        begin
                        left <= data1[1032:1032];
                            middle <= data2[1032:1032];
                            right <= data3[1032:1032];
                        end
                    1033:
                        begin
                        left <= data1[1033:1033];
                            middle <= data2[1033:1033];
                            right <= data3[1033:1033];
                        end
                    1034:
                        begin
                        left <= data1[1034:1034];
                            middle <= data2[1034:1034];
                            right <= data3[1034:1034];
                        end
                    1035:
                        begin
                        left <= data1[1035:1035];
                            middle <= data2[1035:1035];
                            right <= data3[1035:1035];
                        end
                    1036:
                        begin
                        left <= data1[1036:1036];
                            middle <= data2[1036:1036];
                            right <= data3[1036:1036];
                        end
                    1037:
                        begin
                        left <= data1[1037:1037];
                            middle <= data2[1037:1037];
                            right <= data3[1037:1037];
                        end
                    1038:
                        begin
                        left <= data1[1038:1038];
                            middle <= data2[1038:1038];
                            right <= data3[1038:1038];
                        end
                    1039:
                        begin
                        left <= data1[1039:1039];
                            middle <= data2[1039:1039];
                            right <= data3[1039:1039];
                        end
                    1040:
                        begin
                        left <= data1[1040:1040];
                            middle <= data2[1040:1040];
                            right <= data3[1040:1040];
                        end
                    1041:
                        begin
                        left <= data1[1041:1041];
                            middle <= data2[1041:1041];
                            right <= data3[1041:1041];
                        end
                    1042:
                        begin
                        left <= data1[1042:1042];
                            middle <= data2[1042:1042];
                            right <= data3[1042:1042];
                        end
                    1043:
                        begin
                        left <= data1[1043:1043];
                            middle <= data2[1043:1043];
                            right <= data3[1043:1043];
                        end
                    1044:
                        begin
                        left <= data1[1044:1044];
                            middle <= data2[1044:1044];
                            right <= data3[1044:1044];
                        end
                    1045:
                        begin
                        left <= data1[1045:1045];
                            middle <= data2[1045:1045];
                            right <= data3[1045:1045];
                        end
                    1046:
                        begin
                        left <= data1[1046:1046];
                            middle <= data2[1046:1046];
                            right <= data3[1046:1046];
                        end
                    1047:
                        begin
                        left <= data1[1047:1047];
                            middle <= data2[1047:1047];
                            right <= data3[1047:1047];
                        end
                    1048:
                        begin
                        left <= data1[1048:1048];
                            middle <= data2[1048:1048];
                            right <= data3[1048:1048];
                        end
                    1049:
                        begin
                        left <= data1[1049:1049];
                            middle <= data2[1049:1049];
                            right <= data3[1049:1049];
                        end
                    1050:
                        begin
                        left <= data1[1050:1050];
                            middle <= data2[1050:1050];
                            right <= data3[1050:1050];
                        end
                    1051:
                        begin
                        left <= data1[1051:1051];
                            middle <= data2[1051:1051];
                            right <= data3[1051:1051];
                        end
                    1052:
                        begin
                        left <= data1[1052:1052];
                            middle <= data2[1052:1052];
                            right <= data3[1052:1052];
                        end
                    1053:
                        begin
                        left <= data1[1053:1053];
                            middle <= data2[1053:1053];
                            right <= data3[1053:1053];
                        end
                    1054:
                        begin
                        left <= data1[1054:1054];
                            middle <= data2[1054:1054];
                            right <= data3[1054:1054];
                        end
                    1055:
                        begin
                        left <= data1[1055:1055];
                            middle <= data2[1055:1055];
                            right <= data3[1055:1055];
                        end
                    1056:
                        begin
                        left <= data1[1056:1056];
                            middle <= data2[1056:1056];
                            right <= data3[1056:1056];
                        end
                    1057:
                        begin
                        left <= data1[1057:1057];
                            middle <= data2[1057:1057];
                            right <= data3[1057:1057];
                        end
                    1058:
                        begin
                        left <= data1[1058:1058];
                            middle <= data2[1058:1058];
                            right <= data3[1058:1058];
                        end
                    1059:
                        begin
                        left <= data1[1059:1059];
                            middle <= data2[1059:1059];
                            right <= data3[1059:1059];
                        end
                    1060:
                        begin
                        left <= data1[1060:1060];
                            middle <= data2[1060:1060];
                            right <= data3[1060:1060];
                        end
                    1061:
                        begin
                        left <= data1[1061:1061];
                            middle <= data2[1061:1061];
                            right <= data3[1061:1061];
                        end
                    1062:
                        begin
                        left <= data1[1062:1062];
                            middle <= data2[1062:1062];
                            right <= data3[1062:1062];
                        end
                    1063:
                        begin
                        left <= data1[1063:1063];
                            middle <= data2[1063:1063];
                            right <= data3[1063:1063];
                        end
                    1064:
                        begin
                        left <= data1[1064:1064];
                            middle <= data2[1064:1064];
                            right <= data3[1064:1064];
                        end
                    1065:
                        begin
                        left <= data1[1065:1065];
                            middle <= data2[1065:1065];
                            right <= data3[1065:1065];
                        end
                    1066:
                        begin
                        left <= data1[1066:1066];
                            middle <= data2[1066:1066];
                            right <= data3[1066:1066];
                        end
                    1067:
                        begin
                        left <= data1[1067:1067];
                            middle <= data2[1067:1067];
                            right <= data3[1067:1067];
                        end
                    1068:
                        begin
                        left <= data1[1068:1068];
                            middle <= data2[1068:1068];
                            right <= data3[1068:1068];
                        end
                    1069:
                        begin
                        left <= data1[1069:1069];
                            middle <= data2[1069:1069];
                            right <= data3[1069:1069];
                        end
                    1070:
                        begin
                        left <= data1[1070:1070];
                            middle <= data2[1070:1070];
                            right <= data3[1070:1070];
                        end
                    1071:
                        begin
                        left <= data1[1071:1071];
                            middle <= data2[1071:1071];
                            right <= data3[1071:1071];
                        end
                    1072:
                        begin
                        left <= data1[1072:1072];
                            middle <= data2[1072:1072];
                            right <= data3[1072:1072];
                        end
                    1073:
                        begin
                        left <= data1[1073:1073];
                            middle <= data2[1073:1073];
                            right <= data3[1073:1073];
                        end
                    1074:
                        begin
                        left <= data1[1074:1074];
                            middle <= data2[1074:1074];
                            right <= data3[1074:1074];
                        end
                    1075:
                        begin
                        left <= data1[1075:1075];
                            middle <= data2[1075:1075];
                            right <= data3[1075:1075];
                        end
                    1076:
                        begin
                        left <= data1[1076:1076];
                            middle <= data2[1076:1076];
                            right <= data3[1076:1076];
                        end
                    1077:
                        begin
                        left <= data1[1077:1077];
                            middle <= data2[1077:1077];
                            right <= data3[1077:1077];
                        end
                    1078:
                        begin
                        left <= data1[1078:1078];
                            middle <= data2[1078:1078];
                            right <= data3[1078:1078];
                        end
                    1079:
                        begin
                        left <= data1[1079:1079];
                            middle <= data2[1079:1079];
                            right <= data3[1079:1079];
                        end
                    1080:
                        begin
                        left <= data1[1080:1080];
                            middle <= data2[1080:1080];
                            right <= data3[1080:1080];
                        end
                    1081:
                        begin
                        left <= data1[1081:1081];
                            middle <= data2[1081:1081];
                            right <= data3[1081:1081];
                        end
                    1082:
                        begin
                        left <= data1[1082:1082];
                            middle <= data2[1082:1082];
                            right <= data3[1082:1082];
                        end
                    1083:
                        begin
                        left <= data1[1083:1083];
                            middle <= data2[1083:1083];
                            right <= data3[1083:1083];
                        end
                    1084:
                        begin
                        left <= data1[1084:1084];
                            middle <= data2[1084:1084];
                            right <= data3[1084:1084];
                        end
                    1085:
                        begin
                        left <= data1[1085:1085];
                            middle <= data2[1085:1085];
                            right <= data3[1085:1085];
                        end
                    1086:
                        begin
                        left <= data1[1086:1086];
                            middle <= data2[1086:1086];
                            right <= data3[1086:1086];
                        end
                    1087:
                        begin
                        left <= data1[1087:1087];
                            middle <= data2[1087:1087];
                            right <= data3[1087:1087];
                        end
                    1088:
                        begin
                        left <= data1[1088:1088];
                            middle <= data2[1088:1088];
                            right <= data3[1088:1088];
                        end
                    1089:
                        begin
                        left <= data1[1089:1089];
                            middle <= data2[1089:1089];
                            right <= data3[1089:1089];
                        end
                    1090:
                        begin
                        left <= data1[1090:1090];
                            middle <= data2[1090:1090];
                            right <= data3[1090:1090];
                        end
                    1091:
                        begin
                        left <= data1[1091:1091];
                            middle <= data2[1091:1091];
                            right <= data3[1091:1091];
                        end
                    1092:
                        begin
                        left <= data1[1092:1092];
                            middle <= data2[1092:1092];
                            right <= data3[1092:1092];
                        end
                    1093:
                        begin
                        left <= data1[1093:1093];
                            middle <= data2[1093:1093];
                            right <= data3[1093:1093];
                        end
                    1094:
                        begin
                        left <= data1[1094:1094];
                            middle <= data2[1094:1094];
                            right <= data3[1094:1094];
                        end
                    1095:
                        begin
                        left <= data1[1095:1095];
                            middle <= data2[1095:1095];
                            right <= data3[1095:1095];
                        end
                    1096:
                        begin
                        left <= data1[1096:1096];
                            middle <= data2[1096:1096];
                            right <= data3[1096:1096];
                        end
                    1097:
                        begin
                        left <= data1[1097:1097];
                            middle <= data2[1097:1097];
                            right <= data3[1097:1097];
                        end
                    1098:
                        begin
                        left <= data1[1098:1098];
                            middle <= data2[1098:1098];
                            right <= data3[1098:1098];
                        end
                    1099:
                        begin
                        left <= data1[1099:1099];
                            middle <= data2[1099:1099];
                            right <= data3[1099:1099];
                        end
                    1100:
                        begin
                        left <= data1[1100:1100];
                            middle <= data2[1100:1100];
                            right <= data3[1100:1100];
                        end
                    1101:
                        begin
                        left <= data1[1101:1101];
                            middle <= data2[1101:1101];
                            right <= data3[1101:1101];
                        end
                    1102:
                        begin
                        left <= data1[1102:1102];
                            middle <= data2[1102:1102];
                            right <= data3[1102:1102];
                        end
                    1103:
                        begin
                        left <= data1[1103:1103];
                            middle <= data2[1103:1103];
                            right <= data3[1103:1103];
                        end
                    1104:
                        begin
                        left <= data1[1104:1104];
                            middle <= data2[1104:1104];
                            right <= data3[1104:1104];
                        end
                    1105:
                        begin
                        left <= data1[1105:1105];
                            middle <= data2[1105:1105];
                            right <= data3[1105:1105];
                        end
                    1106:
                        begin
                        left <= data1[1106:1106];
                            middle <= data2[1106:1106];
                            right <= data3[1106:1106];
                        end
                    1107:
                        begin
                        left <= data1[1107:1107];
                            middle <= data2[1107:1107];
                            right <= data3[1107:1107];
                        end
                    1108:
                        begin
                        left <= data1[1108:1108];
                            middle <= data2[1108:1108];
                            right <= data3[1108:1108];
                        end
                    1109:
                        begin
                        left <= data1[1109:1109];
                            middle <= data2[1109:1109];
                            right <= data3[1109:1109];
                        end
                    1110:
                        begin
                        left <= data1[1110:1110];
                            middle <= data2[1110:1110];
                            right <= data3[1110:1110];
                        end
                    1111:
                        begin
                        left <= data1[1111:1111];
                            middle <= data2[1111:1111];
                            right <= data3[1111:1111];
                        end
                    1112:
                        begin
                        left <= data1[1112:1112];
                            middle <= data2[1112:1112];
                            right <= data3[1112:1112];
                        end
                    1113:
                        begin
                        left <= data1[1113:1113];
                            middle <= data2[1113:1113];
                            right <= data3[1113:1113];
                        end
                    1114:
                        begin
                        left <= data1[1114:1114];
                            middle <= data2[1114:1114];
                            right <= data3[1114:1114];
                        end
                    1115:
                        begin
                        left <= data1[1115:1115];
                            middle <= data2[1115:1115];
                            right <= data3[1115:1115];
                        end
                    1116:
                        begin
                        left <= data1[1116:1116];
                            middle <= data2[1116:1116];
                            right <= data3[1116:1116];
                        end
                    1117:
                        begin
                        left <= data1[1117:1117];
                            middle <= data2[1117:1117];
                            right <= data3[1117:1117];
                        end
                    1118:
                        begin
                        left <= data1[1118:1118];
                            middle <= data2[1118:1118];
                            right <= data3[1118:1118];
                        end
                    1119:
                        begin
                        left <= data1[1119:1119];
                            middle <= data2[1119:1119];
                            right <= data3[1119:1119];
                        end
                    1120:
                        begin
                        left <= data1[1120:1120];
                            middle <= data2[1120:1120];
                            right <= data3[1120:1120];
                        end
                    1121:
                        begin
                        left <= data1[1121:1121];
                            middle <= data2[1121:1121];
                            right <= data3[1121:1121];
                        end
                    1122:
                        begin
                        left <= data1[1122:1122];
                            middle <= data2[1122:1122];
                            right <= data3[1122:1122];
                        end
                    1123:
                        begin
                        left <= data1[1123:1123];
                            middle <= data2[1123:1123];
                            right <= data3[1123:1123];
                        end
                    1124:
                        begin
                        left <= data1[1124:1124];
                            middle <= data2[1124:1124];
                            right <= data3[1124:1124];
                        end
                    1125:
                        begin
                        left <= data1[1125:1125];
                            middle <= data2[1125:1125];
                            right <= data3[1125:1125];
                        end
                    1126:
                        begin
                        left <= data1[1126:1126];
                            middle <= data2[1126:1126];
                            right <= data3[1126:1126];
                        end
                    1127:
                        begin
                        left <= data1[1127:1127];
                            middle <= data2[1127:1127];
                            right <= data3[1127:1127];
                        end
                    1128:
                        begin
                        left <= data1[1128:1128];
                            middle <= data2[1128:1128];
                            right <= data3[1128:1128];
                        end
                    1129:
                        begin
                        left <= data1[1129:1129];
                            middle <= data2[1129:1129];
                            right <= data3[1129:1129];
                        end
                    1130:
                        begin
                        left <= data1[1130:1130];
                            middle <= data2[1130:1130];
                            right <= data3[1130:1130];
                        end
                    1131:
                        begin
                        left <= data1[1131:1131];
                            middle <= data2[1131:1131];
                            right <= data3[1131:1131];
                        end
                    1132:
                        begin
                        left <= data1[1132:1132];
                            middle <= data2[1132:1132];
                            right <= data3[1132:1132];
                        end
                    1133:
                        begin
                        left <= data1[1133:1133];
                            middle <= data2[1133:1133];
                            right <= data3[1133:1133];
                        end
                    1134:
                        begin
                        left <= data1[1134:1134];
                            middle <= data2[1134:1134];
                            right <= data3[1134:1134];
                        end
                    1135:
                        begin
                        left <= data1[1135:1135];
                            middle <= data2[1135:1135];
                            right <= data3[1135:1135];
                        end
                    1136:
                        begin
                        left <= data1[1136:1136];
                            middle <= data2[1136:1136];
                            right <= data3[1136:1136];
                        end
                    1137:
                        begin
                        left <= data1[1137:1137];
                            middle <= data2[1137:1137];
                            right <= data3[1137:1137];
                        end
                    1138:
                        begin
                        left <= data1[1138:1138];
                            middle <= data2[1138:1138];
                            right <= data3[1138:1138];
                        end
                    1139:
                        begin
                        left <= data1[1139:1139];
                            middle <= data2[1139:1139];
                            right <= data3[1139:1139];
                        end
                    1140:
                        begin
                        left <= data1[1140:1140];
                            middle <= data2[1140:1140];
                            right <= data3[1140:1140];
                        end
                    1141:
                        begin
                        left <= data1[1141:1141];
                            middle <= data2[1141:1141];
                            right <= data3[1141:1141];
                        end
                    1142:
                        begin
                        left <= data1[1142:1142];
                            middle <= data2[1142:1142];
                            right <= data3[1142:1142];
                        end
                    1143:
                        begin
                        left <= data1[1143:1143];
                            middle <= data2[1143:1143];
                            right <= data3[1143:1143];
                        end
                    1144:
                        begin
                        left <= data1[1144:1144];
                            middle <= data2[1144:1144];
                            right <= data3[1144:1144];
                        end
                    1145:
                        begin
                        left <= data1[1145:1145];
                            middle <= data2[1145:1145];
                            right <= data3[1145:1145];
                        end
                    1146:
                        begin
                        left <= data1[1146:1146];
                            middle <= data2[1146:1146];
                            right <= data3[1146:1146];
                        end
                    1147:
                        begin
                        left <= data1[1147:1147];
                            middle <= data2[1147:1147];
                            right <= data3[1147:1147];
                        end
                    1148:
                        begin
                        left <= data1[1148:1148];
                            middle <= data2[1148:1148];
                            right <= data3[1148:1148];
                        end
                    1149:
                        begin
                        left <= data1[1149:1149];
                            middle <= data2[1149:1149];
                            right <= data3[1149:1149];
                        end
                    1150:
                        begin
                        left <= data1[1150:1150];
                            middle <= data2[1150:1150];
                            right <= data3[1150:1150];
                        end
                    1151:
                        begin
                        left <= data1[1151:1151];
                            middle <= data2[1151:1151];
                            right <= data3[1151:1151];
                        end
                    1152:
                        begin
                        left <= data1[1152:1152];
                            middle <= data2[1152:1152];
                            right <= data3[1152:1152];
                        end
                    1153:
                        begin
                        left <= data1[1153:1153];
                            middle <= data2[1153:1153];
                            right <= data3[1153:1153];
                        end
                    1154:
                        begin
                        left <= data1[1154:1154];
                            middle <= data2[1154:1154];
                            right <= data3[1154:1154];
                        end
                    1155:
                        begin
                        left <= data1[1155:1155];
                            middle <= data2[1155:1155];
                            right <= data3[1155:1155];
                        end
                    1156:
                        begin
                        left <= data1[1156:1156];
                            middle <= data2[1156:1156];
                            right <= data3[1156:1156];
                        end
                    1157:
                        begin
                        left <= data1[1157:1157];
                            middle <= data2[1157:1157];
                            right <= data3[1157:1157];
                        end
                    1158:
                        begin
                        left <= data1[1158:1158];
                            middle <= data2[1158:1158];
                            right <= data3[1158:1158];
                        end
                    1159:
                        begin
                        left <= data1[1159:1159];
                            middle <= data2[1159:1159];
                            right <= data3[1159:1159];
                        end
                    1160:
                        begin
                        left <= data1[1160:1160];
                            middle <= data2[1160:1160];
                            right <= data3[1160:1160];
                        end
                    1161:
                        begin
                        left <= data1[1161:1161];
                            middle <= data2[1161:1161];
                            right <= data3[1161:1161];
                        end
                    1162:
                        begin
                        left <= data1[1162:1162];
                            middle <= data2[1162:1162];
                            right <= data3[1162:1162];
                        end
                    1163:
                        begin
                        left <= data1[1163:1163];
                            middle <= data2[1163:1163];
                            right <= data3[1163:1163];
                        end
                    1164:
                        begin
                        left <= data1[1164:1164];
                            middle <= data2[1164:1164];
                            right <= data3[1164:1164];
                        end
                    1165:
                        begin
                        left <= data1[1165:1165];
                            middle <= data2[1165:1165];
                            right <= data3[1165:1165];
                        end
                    1166:
                        begin
                        left <= data1[1166:1166];
                            middle <= data2[1166:1166];
                            right <= data3[1166:1166];
                        end
                    1167:
                        begin
                        left <= data1[1167:1167];
                            middle <= data2[1167:1167];
                            right <= data3[1167:1167];
                        end
                    1168:
                        begin
                        left <= data1[1168:1168];
                            middle <= data2[1168:1168];
                            right <= data3[1168:1168];
                        end
                    1169:
                        begin
                        left <= data1[1169:1169];
                            middle <= data2[1169:1169];
                            right <= data3[1169:1169];
                        end
                    1170:
                        begin
                        left <= data1[1170:1170];
                            middle <= data2[1170:1170];
                            right <= data3[1170:1170];
                        end
                    1171:
                        begin
                        left <= data1[1171:1171];
                            middle <= data2[1171:1171];
                            right <= data3[1171:1171];
                        end
                    1172:
                        begin
                        left <= data1[1172:1172];
                            middle <= data2[1172:1172];
                            right <= data3[1172:1172];
                        end
                    1173:
                        begin
                        left <= data1[1173:1173];
                            middle <= data2[1173:1173];
                            right <= data3[1173:1173];
                        end
                    1174:
                        begin
                        left <= data1[1174:1174];
                            middle <= data2[1174:1174];
                            right <= data3[1174:1174];
                        end
                    1175:
                        begin
                        left <= data1[1175:1175];
                            middle <= data2[1175:1175];
                            right <= data3[1175:1175];
                        end
                    1176:
                        begin
                        left <= data1[1176:1176];
                            middle <= data2[1176:1176];
                            right <= data3[1176:1176];
                        end
                    1177:
                        begin
                        left <= data1[1177:1177];
                            middle <= data2[1177:1177];
                            right <= data3[1177:1177];
                        end
                    1178:
                        begin
                        left <= data1[1178:1178];
                            middle <= data2[1178:1178];
                            right <= data3[1178:1178];
                        end
                    1179:
                        begin
                        left <= data1[1179:1179];
                            middle <= data2[1179:1179];
                            right <= data3[1179:1179];
                        end
                    1180:
                        begin
                        left <= data1[1180:1180];
                            middle <= data2[1180:1180];
                            right <= data3[1180:1180];
                        end
                    1181:
                        begin
                        left <= data1[1181:1181];
                            middle <= data2[1181:1181];
                            right <= data3[1181:1181];
                        end
                    1182:
                        begin
                        left <= data1[1182:1182];
                            middle <= data2[1182:1182];
                            right <= data3[1182:1182];
                        end
                    1183:
                        begin
                        left <= data1[1183:1183];
                            middle <= data2[1183:1183];
                            right <= data3[1183:1183];
                        end
                    1184:
                        begin
                        left <= data1[1184:1184];
                            middle <= data2[1184:1184];
                            right <= data3[1184:1184];
                        end
                    1185:
                        begin
                        left <= data1[1185:1185];
                            middle <= data2[1185:1185];
                            right <= data3[1185:1185];
                        end
                    1186:
                        begin
                        left <= data1[1186:1186];
                            middle <= data2[1186:1186];
                            right <= data3[1186:1186];
                        end
                    1187:
                        begin
                        left <= data1[1187:1187];
                            middle <= data2[1187:1187];
                            right <= data3[1187:1187];
                        end
                    1188:
                        begin
                        left <= data1[1188:1188];
                            middle <= data2[1188:1188];
                            right <= data3[1188:1188];
                        end
                    1189:
                        begin
                        left <= data1[1189:1189];
                            middle <= data2[1189:1189];
                            right <= data3[1189:1189];
                        end
                    1190:
                        begin
                        left <= data1[1190:1190];
                            middle <= data2[1190:1190];
                            right <= data3[1190:1190];
                        end
                    1191:
                        begin
                        left <= data1[1191:1191];
                            middle <= data2[1191:1191];
                            right <= data3[1191:1191];
                        end
                    1192:
                        begin
                        left <= data1[1192:1192];
                            middle <= data2[1192:1192];
                            right <= data3[1192:1192];
                        end
                    1193:
                        begin
                        left <= data1[1193:1193];
                            middle <= data2[1193:1193];
                            right <= data3[1193:1193];
                        end
                    1194:
                        begin
                        left <= data1[1194:1194];
                            middle <= data2[1194:1194];
                            right <= data3[1194:1194];
                        end
                    1195:
                        begin
                        left <= data1[1195:1195];
                            middle <= data2[1195:1195];
                            right <= data3[1195:1195];
                        end
                    1196:
                        begin
                        left <= data1[1196:1196];
                            middle <= data2[1196:1196];
                            right <= data3[1196:1196];
                        end
                    1197:
                        begin
                        left <= data1[1197:1197];
                            middle <= data2[1197:1197];
                            right <= data3[1197:1197];
                        end
                    1198:
                        begin
                        left <= data1[1198:1198];
                            middle <= data2[1198:1198];
                            right <= data3[1198:1198];
                        end
                    1199:
                        begin
                        left <= data1[1199:1199];
                            middle <= data2[1199:1199];
                            right <= data3[1199:1199];
                        end
                    1200:
                        begin
                        left <= data1[1200:1200];
                            middle <= data2[1200:1200];
                            right <= data3[1200:1200];
                        end
                    1201:
                        begin
                        left <= data1[1201:1201];
                            middle <= data2[1201:1201];
                            right <= data3[1201:1201];
                        end
                    1202:
                        begin
                        left <= data1[1202:1202];
                            middle <= data2[1202:1202];
                            right <= data3[1202:1202];
                        end
                    1203:
                        begin
                        left <= data1[1203:1203];
                            middle <= data2[1203:1203];
                            right <= data3[1203:1203];
                        end
                    1204:
                        begin
                        left <= data1[1204:1204];
                            middle <= data2[1204:1204];
                            right <= data3[1204:1204];
                        end
                    1205:
                        begin
                        left <= data1[1205:1205];
                            middle <= data2[1205:1205];
                            right <= data3[1205:1205];
                        end
                    1206:
                        begin
                        left <= data1[1206:1206];
                            middle <= data2[1206:1206];
                            right <= data3[1206:1206];
                        end
                    1207:
                        begin
                        left <= data1[1207:1207];
                            middle <= data2[1207:1207];
                            right <= data3[1207:1207];
                        end
                    1208:
                        begin
                        left <= data1[1208:1208];
                            middle <= data2[1208:1208];
                            right <= data3[1208:1208];
                        end
                    1209:
                        begin
                        left <= data1[1209:1209];
                            middle <= data2[1209:1209];
                            right <= data3[1209:1209];
                        end
                    1210:
                        begin
                        left <= data1[1210:1210];
                            middle <= data2[1210:1210];
                            right <= data3[1210:1210];
                        end
                    1211:
                        begin
                        left <= data1[1211:1211];
                            middle <= data2[1211:1211];
                            right <= data3[1211:1211];
                        end
                    1212:
                        begin
                        left <= data1[1212:1212];
                            middle <= data2[1212:1212];
                            right <= data3[1212:1212];
                        end
                    1213:
                        begin
                        left <= data1[1213:1213];
                            middle <= data2[1213:1213];
                            right <= data3[1213:1213];
                        end
                    1214:
                        begin
                        left <= data1[1214:1214];
                            middle <= data2[1214:1214];
                            right <= data3[1214:1214];
                        end
                    1215:
                        begin
                        left <= data1[1215:1215];
                            middle <= data2[1215:1215];
                            right <= data3[1215:1215];
                        end
                    1216:
                        begin
                        left <= data1[1216:1216];
                            middle <= data2[1216:1216];
                            right <= data3[1216:1216];
                        end
                    1217:
                        begin
                        left <= data1[1217:1217];
                            middle <= data2[1217:1217];
                            right <= data3[1217:1217];
                        end
                    1218:
                        begin
                        left <= data1[1218:1218];
                            middle <= data2[1218:1218];
                            right <= data3[1218:1218];
                        end
                    1219:
                        begin
                        left <= data1[1219:1219];
                            middle <= data2[1219:1219];
                            right <= data3[1219:1219];
                        end
                    1220:
                        begin
                        left <= data1[1220:1220];
                            middle <= data2[1220:1220];
                            right <= data3[1220:1220];
                        end
                    1221:
                        begin
                        left <= data1[1221:1221];
                            middle <= data2[1221:1221];
                            right <= data3[1221:1221];
                        end
                    1222:
                        begin
                        left <= data1[1222:1222];
                            middle <= data2[1222:1222];
                            right <= data3[1222:1222];
                        end
                    1223:
                        begin
                        left <= data1[1223:1223];
                            middle <= data2[1223:1223];
                            right <= data3[1223:1223];
                        end
                    1224:
                        begin
                        left <= data1[1224:1224];
                            middle <= data2[1224:1224];
                            right <= data3[1224:1224];
                        end
                    1225:
                        begin
                        left <= data1[1225:1225];
                            middle <= data2[1225:1225];
                            right <= data3[1225:1225];
                        end
                    1226:
                        begin
                        left <= data1[1226:1226];
                            middle <= data2[1226:1226];
                            right <= data3[1226:1226];
                        end
                    1227:
                        begin
                        left <= data1[1227:1227];
                            middle <= data2[1227:1227];
                            right <= data3[1227:1227];
                        end
                    1228:
                        begin
                        left <= data1[1228:1228];
                            middle <= data2[1228:1228];
                            right <= data3[1228:1228];
                        end
                    1229:
                        begin
                        left <= data1[1229:1229];
                            middle <= data2[1229:1229];
                            right <= data3[1229:1229];
                        end
                    1230:
                        begin
                        left <= data1[1230:1230];
                            middle <= data2[1230:1230];
                            right <= data3[1230:1230];
                        end
                    1231:
                        begin
                        left <= data1[1231:1231];
                            middle <= data2[1231:1231];
                            right <= data3[1231:1231];
                        end
                    1232:
                        begin
                        left <= data1[1232:1232];
                            middle <= data2[1232:1232];
                            right <= data3[1232:1232];
                        end
                    1233:
                        begin
                        left <= data1[1233:1233];
                            middle <= data2[1233:1233];
                            right <= data3[1233:1233];
                        end
                    1234:
                        begin
                        left <= data1[1234:1234];
                            middle <= data2[1234:1234];
                            right <= data3[1234:1234];
                        end
                    1235:
                        begin
                        left <= data1[1235:1235];
                            middle <= data2[1235:1235];
                            right <= data3[1235:1235];
                        end
                    1236:
                        begin
                        left <= data1[1236:1236];
                            middle <= data2[1236:1236];
                            right <= data3[1236:1236];
                        end
                    1237:
                        begin
                        left <= data1[1237:1237];
                            middle <= data2[1237:1237];
                            right <= data3[1237:1237];
                        end
                    1238:
                        begin
                        left <= data1[1238:1238];
                            middle <= data2[1238:1238];
                            right <= data3[1238:1238];
                        end
                    1239:
                        begin
                        left <= data1[1239:1239];
                            middle <= data2[1239:1239];
                            right <= data3[1239:1239];
                        end
                    1240:
                        begin
                        left <= data1[1240:1240];
                            middle <= data2[1240:1240];
                            right <= data3[1240:1240];
                        end
                    1241:
                        begin
                        left <= data1[1241:1241];
                            middle <= data2[1241:1241];
                            right <= data3[1241:1241];
                        end
                    1242:
                        begin
                        left <= data1[1242:1242];
                            middle <= data2[1242:1242];
                            right <= data3[1242:1242];
                        end
                    1243:
                        begin
                        left <= data1[1243:1243];
                            middle <= data2[1243:1243];
                            right <= data3[1243:1243];
                        end
                    1244:
                        begin
                        left <= data1[1244:1244];
                            middle <= data2[1244:1244];
                            right <= data3[1244:1244];
                        end
                    1245:
                        begin
                        left <= data1[1245:1245];
                            middle <= data2[1245:1245];
                            right <= data3[1245:1245];
                        end
                    1246:
                        begin
                        left <= data1[1246:1246];
                            middle <= data2[1246:1246];
                            right <= data3[1246:1246];
                        end
                    1247:
                        begin
                        left <= data1[1247:1247];
                            middle <= data2[1247:1247];
                            right <= data3[1247:1247];
                        end
                    1248:
                        begin
                        left <= data1[1248:1248];
                            middle <= data2[1248:1248];
                            right <= data3[1248:1248];
                        end
                    1249:
                        begin
                        left <= data1[1249:1249];
                            middle <= data2[1249:1249];
                            right <= data3[1249:1249];
                        end
                    1250:
                        begin
                        left <= data1[1250:1250];
                            middle <= data2[1250:1250];
                            right <= data3[1250:1250];
                        end
                    1251:
                        begin
                        left <= data1[1251:1251];
                            middle <= data2[1251:1251];
                            right <= data3[1251:1251];
                        end
                    1252:
                        begin
                        left <= data1[1252:1252];
                            middle <= data2[1252:1252];
                            right <= data3[1252:1252];
                        end
                    1253:
                        begin
                        left <= data1[1253:1253];
                            middle <= data2[1253:1253];
                            right <= data3[1253:1253];
                        end
                    1254:
                        begin
                        left <= data1[1254:1254];
                            middle <= data2[1254:1254];
                            right <= data3[1254:1254];
                        end
                    1255:
                        begin
                        left <= data1[1255:1255];
                            middle <= data2[1255:1255];
                            right <= data3[1255:1255];
                        end
                    1256:
                        begin
                        left <= data1[1256:1256];
                            middle <= data2[1256:1256];
                            right <= data3[1256:1256];
                        end
                    1257:
                        begin
                        left <= data1[1257:1257];
                            middle <= data2[1257:1257];
                            right <= data3[1257:1257];
                        end
                    1258:
                        begin
                        left <= data1[1258:1258];
                            middle <= data2[1258:1258];
                            right <= data3[1258:1258];
                        end
                    1259:
                        begin
                        left <= data1[1259:1259];
                            middle <= data2[1259:1259];
                            right <= data3[1259:1259];
                        end
                    1260:
                        begin
                        left <= data1[1260:1260];
                            middle <= data2[1260:1260];
                            right <= data3[1260:1260];
                        end
                    1261:
                        begin
                        left <= data1[1261:1261];
                            middle <= data2[1261:1261];
                            right <= data3[1261:1261];
                        end
                    1262:
                        begin
                        left <= data1[1262:1262];
                            middle <= data2[1262:1262];
                            right <= data3[1262:1262];
                        end
                    1263:
                        begin
                        left <= data1[1263:1263];
                            middle <= data2[1263:1263];
                            right <= data3[1263:1263];
                        end
                    1264:
                        begin
                        left <= data1[1264:1264];
                            middle <= data2[1264:1264];
                            right <= data3[1264:1264];
                        end
                    1265:
                        begin
                        left <= data1[1265:1265];
                            middle <= data2[1265:1265];
                            right <= data3[1265:1265];
                        end
                    1266:
                        begin
                        left <= data1[1266:1266];
                            middle <= data2[1266:1266];
                            right <= data3[1266:1266];
                        end
                    1267:
                        begin
                        left <= data1[1267:1267];
                            middle <= data2[1267:1267];
                            right <= data3[1267:1267];
                        end
                    1268:
                        begin
                        left <= data1[1268:1268];
                            middle <= data2[1268:1268];
                            right <= data3[1268:1268];
                        end
                    1269:
                        begin
                        left <= data1[1269:1269];
                            middle <= data2[1269:1269];
                            right <= data3[1269:1269];
                        end
                    1270:
                        begin
                        left <= data1[1270:1270];
                            middle <= data2[1270:1270];
                            right <= data3[1270:1270];
                        end
                    1271:
                        begin
                        left <= data1[1271:1271];
                            middle <= data2[1271:1271];
                            right <= data3[1271:1271];
                        end
                    1272:
                        begin
                        left <= data1[1272:1272];
                            middle <= data2[1272:1272];
                            right <= data3[1272:1272];
                        end
                    1273:
                        begin
                        left <= data1[1273:1273];
                            middle <= data2[1273:1273];
                            right <= data3[1273:1273];
                        end
                    1274:
                        begin
                        left <= data1[1274:1274];
                            middle <= data2[1274:1274];
                            right <= data3[1274:1274];
                        end
                    1275:
                        begin
                        left <= data1[1275:1275];
                            middle <= data2[1275:1275];
                            right <= data3[1275:1275];
                        end
                    1276:
                        begin
                        left <= data1[1276:1276];
                            middle <= data2[1276:1276];
                            right <= data3[1276:1276];
                        end
                    1277:
                        begin
                        left <= data1[1277:1277];
                            middle <= data2[1277:1277];
                            right <= data3[1277:1277];
                        end
                    1278:
                        begin
                        left <= data1[1278:1278];
                            middle <= data2[1278:1278];
                            right <= data3[1278:1278];
                        end
                    1279:
                        begin
                        left <= data1[1279:1279];
                            middle <= data2[1279:1279];
                            right <= data3[1279:1279];
                        end
                    1280:
                        begin
                        left <= data1[1280:1280];
                            middle <= data2[1280:1280];
                            right <= data3[1280:1280];
                        end
                    1281:
                        begin
                        left <= data1[1281:1281];
                            middle <= data2[1281:1281];
                            right <= data3[1281:1281];
                        end
                    1282:
                        begin
                        left <= data1[1282:1282];
                            middle <= data2[1282:1282];
                            right <= data3[1282:1282];
                        end
                    1283:
                        begin
                        left <= data1[1283:1283];
                            middle <= data2[1283:1283];
                            right <= data3[1283:1283];
                        end
                    1284:
                        begin
                        left <= data1[1284:1284];
                            middle <= data2[1284:1284];
                            right <= data3[1284:1284];
                        end
                    1285:
                        begin
                        left <= data1[1285:1285];
                            middle <= data2[1285:1285];
                            right <= data3[1285:1285];
                        end
                    1286:
                        begin
                        left <= data1[1286:1286];
                            middle <= data2[1286:1286];
                            right <= data3[1286:1286];
                        end
                    1287:
                        begin
                        left <= data1[1287:1287];
                            middle <= data2[1287:1287];
                            right <= data3[1287:1287];
                        end
                    1288:
                        begin
                        left <= data1[1288:1288];
                            middle <= data2[1288:1288];
                            right <= data3[1288:1288];
                        end
                    1289:
                        begin
                        left <= data1[1289:1289];
                            middle <= data2[1289:1289];
                            right <= data3[1289:1289];
                        end
                    1290:
                        begin
                        left <= data1[1290:1290];
                            middle <= data2[1290:1290];
                            right <= data3[1290:1290];
                        end
                    1291:
                        begin
                        left <= data1[1291:1291];
                            middle <= data2[1291:1291];
                            right <= data3[1291:1291];
                        end
                    1292:
                        begin
                        left <= data1[1292:1292];
                            middle <= data2[1292:1292];
                            right <= data3[1292:1292];
                        end
                    1293:
                        begin
                        left <= data1[1293:1293];
                            middle <= data2[1293:1293];
                            right <= data3[1293:1293];
                        end
                    1294:
                        begin
                        left <= data1[1294:1294];
                            middle <= data2[1294:1294];
                            right <= data3[1294:1294];
                        end
                    1295:
                        begin
                        left <= data1[1295:1295];
                            middle <= data2[1295:1295];
                            right <= data3[1295:1295];
                        end
                    1296:
                        begin
                        left <= data1[1296:1296];
                            middle <= data2[1296:1296];
                            right <= data3[1296:1296];
                        end
                    1297:
                        begin
                        left <= data1[1297:1297];
                            middle <= data2[1297:1297];
                            right <= data3[1297:1297];
                        end
                    1298:
                        begin
                        left <= data1[1298:1298];
                            middle <= data2[1298:1298];
                            right <= data3[1298:1298];
                        end
                    1299:
                        begin
                        left <= data1[1299:1299];
                            middle <= data2[1299:1299];
                            right <= data3[1299:1299];
                        end
                    1300:
                        begin
                        left <= data1[1300:1300];
                            middle <= data2[1300:1300];
                            right <= data3[1300:1300];
                        end
                    1301:
                        begin
                        left <= data1[1301:1301];
                            middle <= data2[1301:1301];
                            right <= data3[1301:1301];
                        end
                    1302:
                        begin
                        left <= data1[1302:1302];
                            middle <= data2[1302:1302];
                            right <= data3[1302:1302];
                        end
                    1303:
                        begin
                        left <= data1[1303:1303];
                            middle <= data2[1303:1303];
                            right <= data3[1303:1303];
                        end
                    1304:
                        begin
                        left <= data1[1304:1304];
                            middle <= data2[1304:1304];
                            right <= data3[1304:1304];
                        end
                    1305:
                        begin
                        left <= data1[1305:1305];
                            middle <= data2[1305:1305];
                            right <= data3[1305:1305];
                        end
                    1306:
                        begin
                        left <= data1[1306:1306];
                            middle <= data2[1306:1306];
                            right <= data3[1306:1306];
                        end
                    1307:
                        begin
                        left <= data1[1307:1307];
                            middle <= data2[1307:1307];
                            right <= data3[1307:1307];
                        end
                    1308:
                        begin
                        left <= data1[1308:1308];
                            middle <= data2[1308:1308];
                            right <= data3[1308:1308];
                        end
                    1309:
                        begin
                        left <= data1[1309:1309];
                            middle <= data2[1309:1309];
                            right <= data3[1309:1309];
                        end
                    1310:
                        begin
                        left <= data1[1310:1310];
                            middle <= data2[1310:1310];
                            right <= data3[1310:1310];
                        end
                    1311:
                        begin
                        left <= data1[1311:1311];
                            middle <= data2[1311:1311];
                            right <= data3[1311:1311];
                        end
                    1312:
                        begin
                        left <= data1[1312:1312];
                            middle <= data2[1312:1312];
                            right <= data3[1312:1312];
                        end
                    1313:
                        begin
                        left <= data1[1313:1313];
                            middle <= data2[1313:1313];
                            right <= data3[1313:1313];
                        end
                    1314:
                        begin
                        left <= data1[1314:1314];
                            middle <= data2[1314:1314];
                            right <= data3[1314:1314];
                        end
                    1315:
                        begin
                        left <= data1[1315:1315];
                            middle <= data2[1315:1315];
                            right <= data3[1315:1315];
                        end
                    1316:
                        begin
                        left <= data1[1316:1316];
                            middle <= data2[1316:1316];
                            right <= data3[1316:1316];
                        end
                    1317:
                        begin
                        left <= data1[1317:1317];
                            middle <= data2[1317:1317];
                            right <= data3[1317:1317];
                        end
                    1318:
                        begin
                        left <= data1[1318:1318];
                            middle <= data2[1318:1318];
                            right <= data3[1318:1318];
                        end
                    1319:
                        begin
                        left <= data1[1319:1319];
                            middle <= data2[1319:1319];
                            right <= data3[1319:1319];
                        end
                    1320:
                        begin
                        left <= data1[1320:1320];
                            middle <= data2[1320:1320];
                            right <= data3[1320:1320];
                        end
                    1321:
                        begin
                        left <= data1[1321:1321];
                            middle <= data2[1321:1321];
                            right <= data3[1321:1321];
                        end
                    1322:
                        begin
                        left <= data1[1322:1322];
                            middle <= data2[1322:1322];
                            right <= data3[1322:1322];
                        end
                    1323:
                        begin
                        left <= data1[1323:1323];
                            middle <= data2[1323:1323];
                            right <= data3[1323:1323];
                        end
                    1324:
                        begin
                        left <= data1[1324:1324];
                            middle <= data2[1324:1324];
                            right <= data3[1324:1324];
                        end
                    1325:
                        begin
                        left <= data1[1325:1325];
                            middle <= data2[1325:1325];
                            right <= data3[1325:1325];
                        end
                    1326:
                        begin
                        left <= data1[1326:1326];
                            middle <= data2[1326:1326];
                            right <= data3[1326:1326];
                        end
                    1327:
                        begin
                        left <= data1[1327:1327];
                            middle <= data2[1327:1327];
                            right <= data3[1327:1327];
                        end
                    1328:
                        begin
                        left <= data1[1328:1328];
                            middle <= data2[1328:1328];
                            right <= data3[1328:1328];
                        end
                    1329:
                        begin
                        left <= data1[1329:1329];
                            middle <= data2[1329:1329];
                            right <= data3[1329:1329];
                        end
                    1330:
                        begin
                        left <= data1[1330:1330];
                            middle <= data2[1330:1330];
                            right <= data3[1330:1330];
                        end
                    1331:
                        begin
                        left <= data1[1331:1331];
                            middle <= data2[1331:1331];
                            right <= data3[1331:1331];
                        end
                    1332:
                        begin
                        left <= data1[1332:1332];
                            middle <= data2[1332:1332];
                            right <= data3[1332:1332];
                        end
                    1333:
                        begin
                        left <= data1[1333:1333];
                            middle <= data2[1333:1333];
                            right <= data3[1333:1333];
                        end
                    1334:
                        begin
                        left <= data1[1334:1334];
                            middle <= data2[1334:1334];
                            right <= data3[1334:1334];
                        end
                    1335:
                        begin
                        left <= data1[1335:1335];
                            middle <= data2[1335:1335];
                            right <= data3[1335:1335];
                        end
                    1336:
                        begin
                        left <= data1[1336:1336];
                            middle <= data2[1336:1336];
                            right <= data3[1336:1336];
                        end
                    1337:
                        begin
                        left <= data1[1337:1337];
                            middle <= data2[1337:1337];
                            right <= data3[1337:1337];
                        end
                    1338:
                        begin
                        left <= data1[1338:1338];
                            middle <= data2[1338:1338];
                            right <= data3[1338:1338];
                        end
                    1339:
                        begin
                        left <= data1[1339:1339];
                            middle <= data2[1339:1339];
                            right <= data3[1339:1339];
                        end
                    1340:
                        begin
                        left <= data1[1340:1340];
                            middle <= data2[1340:1340];
                            right <= data3[1340:1340];
                        end
                    1341:
                        begin
                        left <= data1[1341:1341];
                            middle <= data2[1341:1341];
                            right <= data3[1341:1341];
                        end
                    1342:
                        begin
                        left <= data1[1342:1342];
                            middle <= data2[1342:1342];
                            right <= data3[1342:1342];
                        end
                    1343:
                        begin
                        left <= data1[1343:1343];
                            middle <= data2[1343:1343];
                            right <= data3[1343:1343];
                        end
                    1344:
                        begin
                        left <= data1[1344:1344];
                            middle <= data2[1344:1344];
                            right <= data3[1344:1344];
                        end
                    1345:
                        begin
                        left <= data1[1345:1345];
                            middle <= data2[1345:1345];
                            right <= data3[1345:1345];
                        end
                    1346:
                        begin
                        left <= data1[1346:1346];
                            middle <= data2[1346:1346];
                            right <= data3[1346:1346];
                        end
                    1347:
                        begin
                        left <= data1[1347:1347];
                            middle <= data2[1347:1347];
                            right <= data3[1347:1347];
                        end
                    1348:
                        begin
                        left <= data1[1348:1348];
                            middle <= data2[1348:1348];
                            right <= data3[1348:1348];
                        end
                    1349:
                        begin
                        left <= data1[1349:1349];
                            middle <= data2[1349:1349];
                            right <= data3[1349:1349];
                        end
                    1350:
                        begin
                        left <= data1[1350:1350];
                            middle <= data2[1350:1350];
                            right <= data3[1350:1350];
                        end
                    1351:
                        begin
                        left <= data1[1351:1351];
                            middle <= data2[1351:1351];
                            right <= data3[1351:1351];
                        end
                    1352:
                        begin
                        left <= data1[1352:1352];
                            middle <= data2[1352:1352];
                            right <= data3[1352:1352];
                        end
                    1353:
                        begin
                        left <= data1[1353:1353];
                            middle <= data2[1353:1353];
                            right <= data3[1353:1353];
                        end
                    1354:
                        begin
                        left <= data1[1354:1354];
                            middle <= data2[1354:1354];
                            right <= data3[1354:1354];
                        end
                    1355:
                        begin
                        left <= data1[1355:1355];
                            middle <= data2[1355:1355];
                            right <= data3[1355:1355];
                        end
                    1356:
                        begin
                        left <= data1[1356:1356];
                            middle <= data2[1356:1356];
                            right <= data3[1356:1356];
                        end
                    1357:
                        begin
                        left <= data1[1357:1357];
                            middle <= data2[1357:1357];
                            right <= data3[1357:1357];
                        end
                    1358:
                        begin
                        left <= data1[1358:1358];
                            middle <= data2[1358:1358];
                            right <= data3[1358:1358];
                        end
                    1359:
                        begin
                        left <= data1[1359:1359];
                            middle <= data2[1359:1359];
                            right <= data3[1359:1359];
                        end
                    1360:
                        begin
                        left <= data1[1360:1360];
                            middle <= data2[1360:1360];
                            right <= data3[1360:1360];
                        end
                    1361:
                        begin
                        left <= data1[1361:1361];
                            middle <= data2[1361:1361];
                            right <= data3[1361:1361];
                        end
                    1362:
                        begin
                        left <= data1[1362:1362];
                            middle <= data2[1362:1362];
                            right <= data3[1362:1362];
                        end
                    1363:
                        begin
                        left <= data1[1363:1363];
                            middle <= data2[1363:1363];
                            right <= data3[1363:1363];
                        end
                    1364:
                        begin
                        left <= data1[1364:1364];
                            middle <= data2[1364:1364];
                            right <= data3[1364:1364];
                        end
                    1365:
                        begin
                        left <= data1[1365:1365];
                            middle <= data2[1365:1365];
                            right <= data3[1365:1365];
                        end
                    1366:
                        begin
                        left <= data1[1366:1366];
                            middle <= data2[1366:1366];
                            right <= data3[1366:1366];
                        end
                    1367:
                        begin
                        left <= data1[1367:1367];
                            middle <= data2[1367:1367];
                            right <= data3[1367:1367];
                        end
                    1368:
                        begin
                        left <= data1[1368:1368];
                            middle <= data2[1368:1368];
                            right <= data3[1368:1368];
                        end
                    1369:
                        begin
                        left <= data1[1369:1369];
                            middle <= data2[1369:1369];
                            right <= data3[1369:1369];
                        end
                    1370:
                        begin
                        left <= data1[1370:1370];
                            middle <= data2[1370:1370];
                            right <= data3[1370:1370];
                        end
                    1371:
                        begin
                        left <= data1[1371:1371];
                            middle <= data2[1371:1371];
                            right <= data3[1371:1371];
                        end
                    1372:
                        begin
                        left <= data1[1372:1372];
                            middle <= data2[1372:1372];
                            right <= data3[1372:1372];
                        end
                    1373:
                        begin
                        left <= data1[1373:1373];
                            middle <= data2[1373:1373];
                            right <= data3[1373:1373];
                        end
                    1374:
                        begin
                        left <= data1[1374:1374];
                            middle <= data2[1374:1374];
                            right <= data3[1374:1374];
                        end
                    1375:
                        begin
                        left <= data1[1375:1375];
                            middle <= data2[1375:1375];
                            right <= data3[1375:1375];
                        end
                    1376:
                        begin
                        left <= data1[1376:1376];
                            middle <= data2[1376:1376];
                            right <= data3[1376:1376];
                        end
                    1377:
                        begin
                        left <= data1[1377:1377];
                            middle <= data2[1377:1377];
                            right <= data3[1377:1377];
                        end
                    1378:
                        begin
                        left <= data1[1378:1378];
                            middle <= data2[1378:1378];
                            right <= data3[1378:1378];
                        end
                    1379:
                        begin
                        left <= data1[1379:1379];
                            middle <= data2[1379:1379];
                            right <= data3[1379:1379];
                        end
                    1380:
                        begin
                        left <= data1[1380:1380];
                            middle <= data2[1380:1380];
                            right <= data3[1380:1380];
                        end
                    1381:
                        begin
                        left <= data1[1381:1381];
                            middle <= data2[1381:1381];
                            right <= data3[1381:1381];
                        end
                    1382:
                        begin
                        left <= data1[1382:1382];
                            middle <= data2[1382:1382];
                            right <= data3[1382:1382];
                        end
                    1383:
                        begin
                        left <= data1[1383:1383];
                            middle <= data2[1383:1383];
                            right <= data3[1383:1383];
                        end
                    1384:
                        begin
                        left <= data1[1384:1384];
                            middle <= data2[1384:1384];
                            right <= data3[1384:1384];
                        end
                    1385:
                        begin
                        left <= data1[1385:1385];
                            middle <= data2[1385:1385];
                            right <= data3[1385:1385];
                        end
                    1386:
                        begin
                        left <= data1[1386:1386];
                            middle <= data2[1386:1386];
                            right <= data3[1386:1386];
                        end
                    1387:
                        begin
                        left <= data1[1387:1387];
                            middle <= data2[1387:1387];
                            right <= data3[1387:1387];
                        end
                    1388:
                        begin
                        left <= data1[1388:1388];
                            middle <= data2[1388:1388];
                            right <= data3[1388:1388];
                        end
                    1389:
                        begin
                        left <= data1[1389:1389];
                            middle <= data2[1389:1389];
                            right <= data3[1389:1389];
                        end
                    1390:
                        begin
                        left <= data1[1390:1390];
                            middle <= data2[1390:1390];
                            right <= data3[1390:1390];
                        end
                    1391:
                        begin
                        left <= data1[1391:1391];
                            middle <= data2[1391:1391];
                            right <= data3[1391:1391];
                        end
                    1392:
                        begin
                        left <= data1[1392:1392];
                            middle <= data2[1392:1392];
                            right <= data3[1392:1392];
                        end
                    1393:
                        begin
                        left <= data1[1393:1393];
                            middle <= data2[1393:1393];
                            right <= data3[1393:1393];
                        end
                    1394:
                        begin
                        left <= data1[1394:1394];
                            middle <= data2[1394:1394];
                            right <= data3[1394:1394];
                        end
                    1395:
                        begin
                        left <= data1[1395:1395];
                            middle <= data2[1395:1395];
                            right <= data3[1395:1395];
                        end
                    1396:
                        begin
                        left <= data1[1396:1396];
                            middle <= data2[1396:1396];
                            right <= data3[1396:1396];
                        end
                    1397:
                        begin
                        left <= data1[1397:1397];
                            middle <= data2[1397:1397];
                            right <= data3[1397:1397];
                        end
                    1398:
                        begin
                        left <= data1[1398:1398];
                            middle <= data2[1398:1398];
                            right <= data3[1398:1398];
                        end
                    1399:
                        begin
                        left <= data1[1399:1399];
                            middle <= data2[1399:1399];
                            right <= data3[1399:1399];
                        end
                    1400:
                        begin
                        left <= data1[1400:1400];
                            middle <= data2[1400:1400];
                            right <= data3[1400:1400];
                        end
                    1401:
                        begin
                        left <= data1[1401:1401];
                            middle <= data2[1401:1401];
                            right <= data3[1401:1401];
                        end
                    1402:
                        begin
                        left <= data1[1402:1402];
                            middle <= data2[1402:1402];
                            right <= data3[1402:1402];
                        end
                    1403:
                        begin
                        left <= data1[1403:1403];
                            middle <= data2[1403:1403];
                            right <= data3[1403:1403];
                        end
                    1404:
                        begin
                        left <= data1[1404:1404];
                            middle <= data2[1404:1404];
                            right <= data3[1404:1404];
                        end
                    1405:
                        begin
                        left <= data1[1405:1405];
                            middle <= data2[1405:1405];
                            right <= data3[1405:1405];
                        end
                    1406:
                        begin
                        left <= data1[1406:1406];
                            middle <= data2[1406:1406];
                            right <= data3[1406:1406];
                        end
                    1407:
                        begin
                        left <= data1[1407:1407];
                            middle <= data2[1407:1407];
                            right <= data3[1407:1407];
                        end
                    1408:
                        begin
                        left <= data1[1408:1408];
                            middle <= data2[1408:1408];
                            right <= data3[1408:1408];
                        end
                    1409:
                        begin
                        left <= data1[1409:1409];
                            middle <= data2[1409:1409];
                            right <= data3[1409:1409];
                        end
                    1410:
                        begin
                        left <= data1[1410:1410];
                            middle <= data2[1410:1410];
                            right <= data3[1410:1410];
                        end
                    1411:
                        begin
                        left <= data1[1411:1411];
                            middle <= data2[1411:1411];
                            right <= data3[1411:1411];
                        end
                    1412:
                        begin
                        left <= data1[1412:1412];
                            middle <= data2[1412:1412];
                            right <= data3[1412:1412];
                        end
                    1413:
                        begin
                        left <= data1[1413:1413];
                            middle <= data2[1413:1413];
                            right <= data3[1413:1413];
                        end
                    1414:
                        begin
                        left <= data1[1414:1414];
                            middle <= data2[1414:1414];
                            right <= data3[1414:1414];
                        end
                    1415:
                        begin
                        left <= data1[1415:1415];
                            middle <= data2[1415:1415];
                            right <= data3[1415:1415];
                        end
                    1416:
                        begin
                        left <= data1[1416:1416];
                            middle <= data2[1416:1416];
                            right <= data3[1416:1416];
                        end
                    1417:
                        begin
                        left <= data1[1417:1417];
                            middle <= data2[1417:1417];
                            right <= data3[1417:1417];
                        end
                    1418:
                        begin
                        left <= data1[1418:1418];
                            middle <= data2[1418:1418];
                            right <= data3[1418:1418];
                        end
                    1419:
                        begin
                        left <= data1[1419:1419];
                            middle <= data2[1419:1419];
                            right <= data3[1419:1419];
                        end
                    1420:
                        begin
                        left <= data1[1420:1420];
                            middle <= data2[1420:1420];
                            right <= data3[1420:1420];
                        end
                    1421:
                        begin
                        left <= data1[1421:1421];
                            middle <= data2[1421:1421];
                            right <= data3[1421:1421];
                        end
                    1422:
                        begin
                        left <= data1[1422:1422];
                            middle <= data2[1422:1422];
                            right <= data3[1422:1422];
                        end
                    1423:
                        begin
                        left <= data1[1423:1423];
                            middle <= data2[1423:1423];
                            right <= data3[1423:1423];
                        end
                    1424:
                        begin
                        left <= data1[1424:1424];
                            middle <= data2[1424:1424];
                            right <= data3[1424:1424];
                        end
                    1425:
                        begin
                        left <= data1[1425:1425];
                            middle <= data2[1425:1425];
                            right <= data3[1425:1425];
                        end
                    1426:
                        begin
                        left <= data1[1426:1426];
                            middle <= data2[1426:1426];
                            right <= data3[1426:1426];
                        end
                    1427:
                        begin
                        left <= data1[1427:1427];
                            middle <= data2[1427:1427];
                            right <= data3[1427:1427];
                        end
                    1428:
                        begin
                        left <= data1[1428:1428];
                            middle <= data2[1428:1428];
                            right <= data3[1428:1428];
                        end
                    1429:
                        begin
                        left <= data1[1429:1429];
                            middle <= data2[1429:1429];
                            right <= data3[1429:1429];
                        end
                    1430:
                        begin
                        left <= data1[1430:1430];
                            middle <= data2[1430:1430];
                            right <= data3[1430:1430];
                        end
                    1431:
                        begin
                        left <= data1[1431:1431];
                            middle <= data2[1431:1431];
                            right <= data3[1431:1431];
                        end
                    1432:
                        begin
                        left <= data1[1432:1432];
                            middle <= data2[1432:1432];
                            right <= data3[1432:1432];
                        end
                    1433:
                        begin
                        left <= data1[1433:1433];
                            middle <= data2[1433:1433];
                            right <= data3[1433:1433];
                        end
                    1434:
                        begin
                        left <= data1[1434:1434];
                            middle <= data2[1434:1434];
                            right <= data3[1434:1434];
                        end
                    1435:
                        begin
                        left <= data1[1435:1435];
                            middle <= data2[1435:1435];
                            right <= data3[1435:1435];
                        end
                    1436:
                        begin
                        left <= data1[1436:1436];
                            middle <= data2[1436:1436];
                            right <= data3[1436:1436];
                        end
                    1437:
                        begin
                        left <= data1[1437:1437];
                            middle <= data2[1437:1437];
                            right <= data3[1437:1437];
                        end
                    1438:
                        begin
                        left <= data1[1438:1438];
                            middle <= data2[1438:1438];
                            right <= data3[1438:1438];
                        end
                    1439:
                        begin
                        left <= data1[1439:1439];
                            middle <= data2[1439:1439];
                            right <= data3[1439:1439];
                        end
                    1440:
                        begin
                        left <= data1[1440:1440];
                            middle <= data2[1440:1440];
                            right <= data3[1440:1440];
                        end
                    1441:
                        begin
                        left <= data1[1441:1441];
                            middle <= data2[1441:1441];
                            right <= data3[1441:1441];
                        end
                    1442:
                        begin
                        left <= data1[1442:1442];
                            middle <= data2[1442:1442];
                            right <= data3[1442:1442];
                        end
                    1443:
                        begin
                        left <= data1[1443:1443];
                            middle <= data2[1443:1443];
                            right <= data3[1443:1443];
                        end
                    1444:
                        begin
                        left <= data1[1444:1444];
                            middle <= data2[1444:1444];
                            right <= data3[1444:1444];
                        end
                    1445:
                        begin
                        left <= data1[1445:1445];
                            middle <= data2[1445:1445];
                            right <= data3[1445:1445];
                        end
                    1446:
                        begin
                        left <= data1[1446:1446];
                            middle <= data2[1446:1446];
                            right <= data3[1446:1446];
                        end
                    1447:
                        begin
                        left <= data1[1447:1447];
                            middle <= data2[1447:1447];
                            right <= data3[1447:1447];
                        end
                    1448:
                        begin
                        left <= data1[1448:1448];
                            middle <= data2[1448:1448];
                            right <= data3[1448:1448];
                        end
                    1449:
                        begin
                        left <= data1[1449:1449];
                            middle <= data2[1449:1449];
                            right <= data3[1449:1449];
                        end
                    1450:
                        begin
                        left <= data1[1450:1450];
                            middle <= data2[1450:1450];
                            right <= data3[1450:1450];
                        end
                    1451:
                        begin
                        left <= data1[1451:1451];
                            middle <= data2[1451:1451];
                            right <= data3[1451:1451];
                        end
                    1452:
                        begin
                        left <= data1[1452:1452];
                            middle <= data2[1452:1452];
                            right <= data3[1452:1452];
                        end
                    1453:
                        begin
                        left <= data1[1453:1453];
                            middle <= data2[1453:1453];
                            right <= data3[1453:1453];
                        end
                    1454:
                        begin
                        left <= data1[1454:1454];
                            middle <= data2[1454:1454];
                            right <= data3[1454:1454];
                        end
                    1455:
                        begin
                        left <= data1[1455:1455];
                            middle <= data2[1455:1455];
                            right <= data3[1455:1455];
                        end
                    1456:
                        begin
                        left <= data1[1456:1456];
                            middle <= data2[1456:1456];
                            right <= data3[1456:1456];
                        end
                    1457:
                        begin
                        left <= data1[1457:1457];
                            middle <= data2[1457:1457];
                            right <= data3[1457:1457];
                        end
                    1458:
                        begin
                        left <= data1[1458:1458];
                            middle <= data2[1458:1458];
                            right <= data3[1458:1458];
                        end
                    1459:
                        begin
                        left <= data1[1459:1459];
                            middle <= data2[1459:1459];
                            right <= data3[1459:1459];
                        end
                    1460:
                        begin
                        left <= data1[1460:1460];
                            middle <= data2[1460:1460];
                            right <= data3[1460:1460];
                        end
                    1461:
                        begin
                        left <= data1[1461:1461];
                            middle <= data2[1461:1461];
                            right <= data3[1461:1461];
                        end
                    1462:
                        begin
                        left <= data1[1462:1462];
                            middle <= data2[1462:1462];
                            right <= data3[1462:1462];
                        end
                    1463:
                        begin
                        left <= data1[1463:1463];
                            middle <= data2[1463:1463];
                            right <= data3[1463:1463];
                        end
                    1464:
                        begin
                        left <= data1[1464:1464];
                            middle <= data2[1464:1464];
                            right <= data3[1464:1464];
                        end
                    1465:
                        begin
                        left <= data1[1465:1465];
                            middle <= data2[1465:1465];
                            right <= data3[1465:1465];
                        end
                    1466:
                        begin
                        left <= data1[1466:1466];
                            middle <= data2[1466:1466];
                            right <= data3[1466:1466];
                        end
                    1467:
                        begin
                        left <= data1[1467:1467];
                            middle <= data2[1467:1467];
                            right <= data3[1467:1467];
                        end
                    1468:
                        begin
                        left <= data1[1468:1468];
                            middle <= data2[1468:1468];
                            right <= data3[1468:1468];
                        end
                    1469:
                        begin
                        left <= data1[1469:1469];
                            middle <= data2[1469:1469];
                            right <= data3[1469:1469];
                        end
                    1470:
                        begin
                        left <= data1[1470:1470];
                            middle <= data2[1470:1470];
                            right <= data3[1470:1470];
                        end
                    1471:
                        begin
                        left <= data1[1471:1471];
                            middle <= data2[1471:1471];
                            right <= data3[1471:1471];
                        end
                    1472:
                        begin
                        left <= data1[1472:1472];
                            middle <= data2[1472:1472];
                            right <= data3[1472:1472];
                        end
                    1473:
                        begin
                        left <= data1[1473:1473];
                            middle <= data2[1473:1473];
                            right <= data3[1473:1473];
                        end
                    1474:
                        begin
                        left <= data1[1474:1474];
                            middle <= data2[1474:1474];
                            right <= data3[1474:1474];
                        end
                    1475:
                        begin
                        left <= data1[1475:1475];
                            middle <= data2[1475:1475];
                            right <= data3[1475:1475];
                        end
                    1476:
                        begin
                        left <= data1[1476:1476];
                            middle <= data2[1476:1476];
                            right <= data3[1476:1476];
                        end
                    1477:
                        begin
                        left <= data1[1477:1477];
                            middle <= data2[1477:1477];
                            right <= data3[1477:1477];
                        end
                    1478:
                        begin
                        left <= data1[1478:1478];
                            middle <= data2[1478:1478];
                            right <= data3[1478:1478];
                        end
                    1479:
                        begin
                        left <= data1[1479:1479];
                            middle <= data2[1479:1479];
                            right <= data3[1479:1479];
                        end
                    1480:
                        begin
                        left <= data1[1480:1480];
                            middle <= data2[1480:1480];
                            right <= data3[1480:1480];
                        end
                    1481:
                        begin
                        left <= data1[1481:1481];
                            middle <= data2[1481:1481];
                            right <= data3[1481:1481];
                        end
                    1482:
                        begin
                        left <= data1[1482:1482];
                            middle <= data2[1482:1482];
                            right <= data3[1482:1482];
                        end
                    1483:
                        begin
                        left <= data1[1483:1483];
                            middle <= data2[1483:1483];
                            right <= data3[1483:1483];
                        end
                    1484:
                        begin
                        left <= data1[1484:1484];
                            middle <= data2[1484:1484];
                            right <= data3[1484:1484];
                        end
                    1485:
                        begin
                        left <= data1[1485:1485];
                            middle <= data2[1485:1485];
                            right <= data3[1485:1485];
                        end
                    1486:
                        begin
                        left <= data1[1486:1486];
                            middle <= data2[1486:1486];
                            right <= data3[1486:1486];
                        end
                    1487:
                        begin
                        left <= data1[1487:1487];
                            middle <= data2[1487:1487];
                            right <= data3[1487:1487];
                        end
                    1488:
                        begin
                        left <= data1[1488:1488];
                            middle <= data2[1488:1488];
                            right <= data3[1488:1488];
                        end
                    1489:
                        begin
                        left <= data1[1489:1489];
                            middle <= data2[1489:1489];
                            right <= data3[1489:1489];
                        end
                    1490:
                        begin
                        left <= data1[1490:1490];
                            middle <= data2[1490:1490];
                            right <= data3[1490:1490];
                        end
                    1491:
                        begin
                        left <= data1[1491:1491];
                            middle <= data2[1491:1491];
                            right <= data3[1491:1491];
                        end
                    1492:
                        begin
                        left <= data1[1492:1492];
                            middle <= data2[1492:1492];
                            right <= data3[1492:1492];
                        end
                    1493:
                        begin
                        left <= data1[1493:1493];
                            middle <= data2[1493:1493];
                            right <= data3[1493:1493];
                        end
                    1494:
                        begin
                        left <= data1[1494:1494];
                            middle <= data2[1494:1494];
                            right <= data3[1494:1494];
                        end
                    1495:
                        begin
                        left <= data1[1495:1495];
                            middle <= data2[1495:1495];
                            right <= data3[1495:1495];
                        end
                    1496:
                        begin
                        left <= data1[1496:1496];
                            middle <= data2[1496:1496];
                            right <= data3[1496:1496];
                        end
                    1497:
                        begin
                        left <= data1[1497:1497];
                            middle <= data2[1497:1497];
                            right <= data3[1497:1497];
                        end
                    1498:
                        begin
                        left <= data1[1498:1498];
                            middle <= data2[1498:1498];
                            right <= data3[1498:1498];
                        end
                    1499:
                        begin
                        left <= data1[1499:1499];
                            middle <= data2[1499:1499];
                            right <= data3[1499:1499];
                        end
                    1500:
                        begin
                        left <= data1[1500:1500];
                            middle <= data2[1500:1500];
                            right <= data3[1500:1500];
                        end
                    1501:
                        begin
                        left <= data1[1501:1501];
                            middle <= data2[1501:1501];
                            right <= data3[1501:1501];
                        end
                    1502:
                        begin
                        left <= data1[1502:1502];
                            middle <= data2[1502:1502];
                            right <= data3[1502:1502];
                        end
                    1503:
                        begin
                        left <= data1[1503:1503];
                            middle <= data2[1503:1503];
                            right <= data3[1503:1503];
                        end
                    1504:
                        begin
                        left <= data1[1504:1504];
                            middle <= data2[1504:1504];
                            right <= data3[1504:1504];
                        end
                    1505:
                        begin
                        left <= data1[1505:1505];
                            middle <= data2[1505:1505];
                            right <= data3[1505:1505];
                        end
                    1506:
                        begin
                        left <= data1[1506:1506];
                            middle <= data2[1506:1506];
                            right <= data3[1506:1506];
                        end
                    1507:
                        begin
                        left <= data1[1507:1507];
                            middle <= data2[1507:1507];
                            right <= data3[1507:1507];
                        end
                    1508:
                        begin
                        left <= data1[1508:1508];
                            middle <= data2[1508:1508];
                            right <= data3[1508:1508];
                        end
                    1509:
                        begin
                        left <= data1[1509:1509];
                            middle <= data2[1509:1509];
                            right <= data3[1509:1509];
                        end
                    1510:
                        begin
                        left <= data1[1510:1510];
                            middle <= data2[1510:1510];
                            right <= data3[1510:1510];
                        end
                    1511:
                        begin
                        left <= data1[1511:1511];
                            middle <= data2[1511:1511];
                            right <= data3[1511:1511];
                        end
                    1512:
                        begin
                        left <= data1[1512:1512];
                            middle <= data2[1512:1512];
                            right <= data3[1512:1512];
                        end
                    1513:
                        begin
                        left <= data1[1513:1513];
                            middle <= data2[1513:1513];
                            right <= data3[1513:1513];
                        end
                    1514:
                        begin
                        left <= data1[1514:1514];
                            middle <= data2[1514:1514];
                            right <= data3[1514:1514];
                        end
                    1515:
                        begin
                        left <= data1[1515:1515];
                            middle <= data2[1515:1515];
                            right <= data3[1515:1515];
                        end
                    1516:
                        begin
                        left <= data1[1516:1516];
                            middle <= data2[1516:1516];
                            right <= data3[1516:1516];
                        end
                    1517:
                        begin
                        left <= data1[1517:1517];
                            middle <= data2[1517:1517];
                            right <= data3[1517:1517];
                        end
                    1518:
                        begin
                        left <= data1[1518:1518];
                            middle <= data2[1518:1518];
                            right <= data3[1518:1518];
                        end
                    1519:
                        begin
                        left <= data1[1519:1519];
                            middle <= data2[1519:1519];
                            right <= data3[1519:1519];
                        end
                    1520:
                        begin
                        left <= data1[1520:1520];
                            middle <= data2[1520:1520];
                            right <= data3[1520:1520];
                        end
                    1521:
                        begin
                        left <= data1[1521:1521];
                            middle <= data2[1521:1521];
                            right <= data3[1521:1521];
                        end
                    1522:
                        begin
                        left <= data1[1522:1522];
                            middle <= data2[1522:1522];
                            right <= data3[1522:1522];
                        end
                    1523:
                        begin
                        left <= data1[1523:1523];
                            middle <= data2[1523:1523];
                            right <= data3[1523:1523];
                        end
                    1524:
                        begin
                        left <= data1[1524:1524];
                            middle <= data2[1524:1524];
                            right <= data3[1524:1524];
                        end
                    1525:
                        begin
                        left <= data1[1525:1525];
                            middle <= data2[1525:1525];
                            right <= data3[1525:1525];
                        end
                    1526:
                        begin
                        left <= data1[1526:1526];
                            middle <= data2[1526:1526];
                            right <= data3[1526:1526];
                        end
                    1527:
                        begin
                        left <= data1[1527:1527];
                            middle <= data2[1527:1527];
                            right <= data3[1527:1527];
                        end
                    1528:
                        begin
                        left <= data1[1528:1528];
                            middle <= data2[1528:1528];
                            right <= data3[1528:1528];
                        end
                    1529:
                        begin
                        left <= data1[1529:1529];
                            middle <= data2[1529:1529];
                            right <= data3[1529:1529];
                        end
                    1530:
                        begin
                        left <= data1[1530:1530];
                            middle <= data2[1530:1530];
                            right <= data3[1530:1530];
                        end
                    1531:
                        begin
                        left <= data1[1531:1531];
                            middle <= data2[1531:1531];
                            right <= data3[1531:1531];
                        end
                    1532:
                        begin
                        left <= data1[1532:1532];
                            middle <= data2[1532:1532];
                            right <= data3[1532:1532];
                        end
                    1533:
                        begin
                        left <= data1[1533:1533];
                            middle <= data2[1533:1533];
                            right <= data3[1533:1533];
                        end
                    1534:
                        begin
                        left <= data1[1534:1534];
                            middle <= data2[1534:1534];
                            right <= data3[1534:1534];
                        end
                    1535:
                        begin
                        left <= data1[1535:1535];
                            middle <= data2[1535:1535];
                            right <= data3[1535:1535];
                        end
                    1536:
                        begin
                        left <= data1[1536:1536];
                            middle <= data2[1536:1536];
                            right <= data3[1536:1536];
                        end
                    1537:
                        begin
                        left <= data1[1537:1537];
                            middle <= data2[1537:1537];
                            right <= data3[1537:1537];
                        end
                    1538:
                        begin
                        left <= data1[1538:1538];
                            middle <= data2[1538:1538];
                            right <= data3[1538:1538];
                        end
                    1539:
                        begin
                        left <= data1[1539:1539];
                            middle <= data2[1539:1539];
                            right <= data3[1539:1539];
                        end
                    1540:
                        begin
                        left <= data1[1540:1540];
                            middle <= data2[1540:1540];
                            right <= data3[1540:1540];
                        end
                    1541:
                        begin
                        left <= data1[1541:1541];
                            middle <= data2[1541:1541];
                            right <= data3[1541:1541];
                        end
                    1542:
                        begin
                        left <= data1[1542:1542];
                            middle <= data2[1542:1542];
                            right <= data3[1542:1542];
                        end
                    1543:
                        begin
                        left <= data1[1543:1543];
                            middle <= data2[1543:1543];
                            right <= data3[1543:1543];
                        end
                    1544:
                        begin
                        left <= data1[1544:1544];
                            middle <= data2[1544:1544];
                            right <= data3[1544:1544];
                        end
                    1545:
                        begin
                        left <= data1[1545:1545];
                            middle <= data2[1545:1545];
                            right <= data3[1545:1545];
                        end
                    1546:
                        begin
                        left <= data1[1546:1546];
                            middle <= data2[1546:1546];
                            right <= data3[1546:1546];
                        end
                    1547:
                        begin
                        left <= data1[1547:1547];
                            middle <= data2[1547:1547];
                            right <= data3[1547:1547];
                        end
                    1548:
                        begin
                        left <= data1[1548:1548];
                            middle <= data2[1548:1548];
                            right <= data3[1548:1548];
                        end
                    1549:
                        begin
                        left <= data1[1549:1549];
                            middle <= data2[1549:1549];
                            right <= data3[1549:1549];
                        end
                    1550:
                        begin
                        left <= data1[1550:1550];
                            middle <= data2[1550:1550];
                            right <= data3[1550:1550];
                        end
                    1551:
                        begin
                        left <= data1[1551:1551];
                            middle <= data2[1551:1551];
                            right <= data3[1551:1551];
                        end
                    1552:
                        begin
                        left <= data1[1552:1552];
                            middle <= data2[1552:1552];
                            right <= data3[1552:1552];
                        end
                    1553:
                        begin
                        left <= data1[1553:1553];
                            middle <= data2[1553:1553];
                            right <= data3[1553:1553];
                        end
                    1554:
                        begin
                        left <= data1[1554:1554];
                            middle <= data2[1554:1554];
                            right <= data3[1554:1554];
                        end
                    1555:
                        begin
                        left <= data1[1555:1555];
                            middle <= data2[1555:1555];
                            right <= data3[1555:1555];
                        end
                    1556:
                        begin
                        left <= data1[1556:1556];
                            middle <= data2[1556:1556];
                            right <= data3[1556:1556];
                        end
                    1557:
                        begin
                        left <= data1[1557:1557];
                            middle <= data2[1557:1557];
                            right <= data3[1557:1557];
                        end
                    1558:
                        begin
                        left <= data1[1558:1558];
                            middle <= data2[1558:1558];
                            right <= data3[1558:1558];
                        end
                    1559:
                        begin
                        left <= data1[1559:1559];
                            middle <= data2[1559:1559];
                            right <= data3[1559:1559];
                        end
                    1560:
                        begin
                        left <= data1[1560:1560];
                            middle <= data2[1560:1560];
                            right <= data3[1560:1560];
                        end
                    1561:
                        begin
                        left <= data1[1561:1561];
                            middle <= data2[1561:1561];
                            right <= data3[1561:1561];
                        end
                    1562:
                        begin
                        left <= data1[1562:1562];
                            middle <= data2[1562:1562];
                            right <= data3[1562:1562];
                        end
                    1563:
                        begin
                        left <= data1[1563:1563];
                            middle <= data2[1563:1563];
                            right <= data3[1563:1563];
                        end
                    1564:
                        begin
                        left <= data1[1564:1564];
                            middle <= data2[1564:1564];
                            right <= data3[1564:1564];
                        end
                    1565:
                        begin
                        left <= data1[1565:1565];
                            middle <= data2[1565:1565];
                            right <= data3[1565:1565];
                        end
                    1566:
                        begin
                        left <= data1[1566:1566];
                            middle <= data2[1566:1566];
                            right <= data3[1566:1566];
                        end
                    1567:
                        begin
                        left <= data1[1567:1567];
                            middle <= data2[1567:1567];
                            right <= data3[1567:1567];
                        end
                    1568:
                        begin
                        left <= data1[1568:1568];
                            middle <= data2[1568:1568];
                            right <= data3[1568:1568];
                        end
                    1569:
                        begin
                        left <= data1[1569:1569];
                            middle <= data2[1569:1569];
                            right <= data3[1569:1569];
                        end
                    1570:
                        begin
                        left <= data1[1570:1570];
                            middle <= data2[1570:1570];
                            right <= data3[1570:1570];
                        end
                    1571:
                        begin
                        left <= data1[1571:1571];
                            middle <= data2[1571:1571];
                            right <= data3[1571:1571];
                        end
                    1572:
                        begin
                        left <= data1[1572:1572];
                            middle <= data2[1572:1572];
                            right <= data3[1572:1572];
                        end
                    1573:
                        begin
                        left <= data1[1573:1573];
                            middle <= data2[1573:1573];
                            right <= data3[1573:1573];
                        end
                    1574:
                        begin
                        left <= data1[1574:1574];
                            middle <= data2[1574:1574];
                            right <= data3[1574:1574];
                        end
                    1575:
                        begin
                        left <= data1[1575:1575];
                            middle <= data2[1575:1575];
                            right <= data3[1575:1575];
                        end
                    1576:
                        begin
                        left <= data1[1576:1576];
                            middle <= data2[1576:1576];
                            right <= data3[1576:1576];
                        end
                    1577:
                        begin
                        left <= data1[1577:1577];
                            middle <= data2[1577:1577];
                            right <= data3[1577:1577];
                        end
                    1578:
                        begin
                        left <= data1[1578:1578];
                            middle <= data2[1578:1578];
                            right <= data3[1578:1578];
                        end
                    1579:
                        begin
                        left <= data1[1579:1579];
                            middle <= data2[1579:1579];
                            right <= data3[1579:1579];
                        end
                    1580:
                        begin
                        left <= data1[1580:1580];
                            middle <= data2[1580:1580];
                            right <= data3[1580:1580];
                        end
                    1581:
                        begin
                        left <= data1[1581:1581];
                            middle <= data2[1581:1581];
                            right <= data3[1581:1581];
                        end
                    1582:
                        begin
                        left <= data1[1582:1582];
                            middle <= data2[1582:1582];
                            right <= data3[1582:1582];
                        end
                    1583:
                        begin
                        left <= data1[1583:1583];
                            middle <= data2[1583:1583];
                            right <= data3[1583:1583];
                        end
                    1584:
                        begin
                        left <= data1[1584:1584];
                            middle <= data2[1584:1584];
                            right <= data3[1584:1584];
                        end
                    1585:
                        begin
                        left <= data1[1585:1585];
                            middle <= data2[1585:1585];
                            right <= data3[1585:1585];
                        end
                    1586:
                        begin
                        left <= data1[1586:1586];
                            middle <= data2[1586:1586];
                            right <= data3[1586:1586];
                        end
                    1587:
                        begin
                        left <= data1[1587:1587];
                            middle <= data2[1587:1587];
                            right <= data3[1587:1587];
                        end
                    1588:
                        begin
                        left <= data1[1588:1588];
                            middle <= data2[1588:1588];
                            right <= data3[1588:1588];
                        end
                    1589:
                        begin
                        left <= data1[1589:1589];
                            middle <= data2[1589:1589];
                            right <= data3[1589:1589];
                        end
                    1590:
                        begin
                        left <= data1[1590:1590];
                            middle <= data2[1590:1590];
                            right <= data3[1590:1590];
                        end
                    1591:
                        begin
                        left <= data1[1591:1591];
                            middle <= data2[1591:1591];
                            right <= data3[1591:1591];
                        end
                    1592:
                        begin
                        left <= data1[1592:1592];
                            middle <= data2[1592:1592];
                            right <= data3[1592:1592];
                        end
                    1593:
                        begin
                        left <= data1[1593:1593];
                            middle <= data2[1593:1593];
                            right <= data3[1593:1593];
                        end
                    1594:
                        begin
                        left <= data1[1594:1594];
                            middle <= data2[1594:1594];
                            right <= data3[1594:1594];
                        end
                    1595:
                        begin
                        left <= data1[1595:1595];
                            middle <= data2[1595:1595];
                            right <= data3[1595:1595];
                        end
                    1596:
                        begin
                        left <= data1[1596:1596];
                            middle <= data2[1596:1596];
                            right <= data3[1596:1596];
                        end
                    1597:
                        begin
                        left <= data1[1597:1597];
                            middle <= data2[1597:1597];
                            right <= data3[1597:1597];
                        end
                    1598:
                        begin
                        left <= data1[1598:1598];
                            middle <= data2[1598:1598];
                            right <= data3[1598:1598];
                        end
                    1599:
                        begin
                        left <= data1[1599:1599];
                            middle <= data2[1599:1599];
                            right <= data3[1599:1599];
                        end
                    1600:
                        begin
                        left <= data1[1600:1600];
                            middle <= data2[1600:1600];
                            right <= data3[1600:1600];
                        end
                    1601:
                        begin
                        left <= data1[1601:1601];
                            middle <= data2[1601:1601];
                            right <= data3[1601:1601];
                        end
                    1602:
                        begin
                        left <= data1[1602:1602];
                            middle <= data2[1602:1602];
                            right <= data3[1602:1602];
                        end
                    1603:
                        begin
                        left <= data1[1603:1603];
                            middle <= data2[1603:1603];
                            right <= data3[1603:1603];
                        end
                    1604:
                        begin
                        left <= data1[1604:1604];
                            middle <= data2[1604:1604];
                            right <= data3[1604:1604];
                        end
                    1605:
                        begin
                        left <= data1[1605:1605];
                            middle <= data2[1605:1605];
                            right <= data3[1605:1605];
                        end
                    1606:
                        begin
                        left <= data1[1606:1606];
                            middle <= data2[1606:1606];
                            right <= data3[1606:1606];
                        end
                    1607:
                        begin
                        left <= data1[1607:1607];
                            middle <= data2[1607:1607];
                            right <= data3[1607:1607];
                        end
                    1608:
                        begin
                        left <= data1[1608:1608];
                            middle <= data2[1608:1608];
                            right <= data3[1608:1608];
                        end
                    1609:
                        begin
                        left <= data1[1609:1609];
                            middle <= data2[1609:1609];
                            right <= data3[1609:1609];
                        end
                    1610:
                        begin
                        left <= data1[1610:1610];
                            middle <= data2[1610:1610];
                            right <= data3[1610:1610];
                        end
                    1611:
                        begin
                        left <= data1[1611:1611];
                            middle <= data2[1611:1611];
                            right <= data3[1611:1611];
                        end
                    1612:
                        begin
                        left <= data1[1612:1612];
                            middle <= data2[1612:1612];
                            right <= data3[1612:1612];
                        end
                    1613:
                        begin
                        left <= data1[1613:1613];
                            middle <= data2[1613:1613];
                            right <= data3[1613:1613];
                        end
                    1614:
                        begin
                        left <= data1[1614:1614];
                            middle <= data2[1614:1614];
                            right <= data3[1614:1614];
                        end
                    1615:
                        begin
                        left <= data1[1615:1615];
                            middle <= data2[1615:1615];
                            right <= data3[1615:1615];
                        end
                    1616:
                        begin
                        left <= data1[1616:1616];
                            middle <= data2[1616:1616];
                            right <= data3[1616:1616];
                        end
                    1617:
                        begin
                        left <= data1[1617:1617];
                            middle <= data2[1617:1617];
                            right <= data3[1617:1617];
                        end
                    1618:
                        begin
                        left <= data1[1618:1618];
                            middle <= data2[1618:1618];
                            right <= data3[1618:1618];
                        end
                    1619:
                        begin
                        left <= data1[1619:1619];
                            middle <= data2[1619:1619];
                            right <= data3[1619:1619];
                        end
                    1620:
                        begin
                        left <= data1[1620:1620];
                            middle <= data2[1620:1620];
                            right <= data3[1620:1620];
                        end
                    1621:
                        begin
                        left <= data1[1621:1621];
                            middle <= data2[1621:1621];
                            right <= data3[1621:1621];
                        end
                    1622:
                        begin
                        left <= data1[1622:1622];
                            middle <= data2[1622:1622];
                            right <= data3[1622:1622];
                        end
                    1623:
                        begin
                        left <= data1[1623:1623];
                            middle <= data2[1623:1623];
                            right <= data3[1623:1623];
                        end
                    1624:
                        begin
                        left <= data1[1624:1624];
                            middle <= data2[1624:1624];
                            right <= data3[1624:1624];
                        end
                    1625:
                        begin
                        left <= data1[1625:1625];
                            middle <= data2[1625:1625];
                            right <= data3[1625:1625];
                        end
                    1626:
                        begin
                        left <= data1[1626:1626];
                            middle <= data2[1626:1626];
                            right <= data3[1626:1626];
                        end
                    1627:
                        begin
                        left <= data1[1627:1627];
                            middle <= data2[1627:1627];
                            right <= data3[1627:1627];
                        end
                    1628:
                        begin
                        left <= data1[1628:1628];
                            middle <= data2[1628:1628];
                            right <= data3[1628:1628];
                        end
                    1629:
                        begin
                        left <= data1[1629:1629];
                            middle <= data2[1629:1629];
                            right <= data3[1629:1629];
                        end
                    1630:
                        begin
                        left <= data1[1630:1630];
                            middle <= data2[1630:1630];
                            right <= data3[1630:1630];
                        end
                    1631:
                        begin
                        left <= data1[1631:1631];
                            middle <= data2[1631:1631];
                            right <= data3[1631:1631];
                        end
                    1632:
                        begin
                        left <= data1[1632:1632];
                            middle <= data2[1632:1632];
                            right <= data3[1632:1632];
                        end
                    1633:
                        begin
                        left <= data1[1633:1633];
                            middle <= data2[1633:1633];
                            right <= data3[1633:1633];
                        end
                    1634:
                        begin
                        left <= data1[1634:1634];
                            middle <= data2[1634:1634];
                            right <= data3[1634:1634];
                        end
                    1635:
                        begin
                        left <= data1[1635:1635];
                            middle <= data2[1635:1635];
                            right <= data3[1635:1635];
                        end
                    1636:
                        begin
                        left <= data1[1636:1636];
                            middle <= data2[1636:1636];
                            right <= data3[1636:1636];
                        end
                    1637:
                        begin
                        left <= data1[1637:1637];
                            middle <= data2[1637:1637];
                            right <= data3[1637:1637];
                        end
                    1638:
                        begin
                        left <= data1[1638:1638];
                            middle <= data2[1638:1638];
                            right <= data3[1638:1638];
                        end
                    1639:
                        begin
                        left <= data1[1639:1639];
                            middle <= data2[1639:1639];
                            right <= data3[1639:1639];
                        end
                    1640:
                        begin
                        left <= data1[1640:1640];
                            middle <= data2[1640:1640];
                            right <= data3[1640:1640];
                        end
                    1641:
                        begin
                        left <= data1[1641:1641];
                            middle <= data2[1641:1641];
                            right <= data3[1641:1641];
                        end
                    1642:
                        begin
                        left <= data1[1642:1642];
                            middle <= data2[1642:1642];
                            right <= data3[1642:1642];
                        end
                    1643:
                        begin
                        left <= data1[1643:1643];
                            middle <= data2[1643:1643];
                            right <= data3[1643:1643];
                        end
                    1644:
                        begin
                        left <= data1[1644:1644];
                            middle <= data2[1644:1644];
                            right <= data3[1644:1644];
                        end
                    1645:
                        begin
                        left <= data1[1645:1645];
                            middle <= data2[1645:1645];
                            right <= data3[1645:1645];
                        end
                    1646:
                        begin
                        left <= data1[1646:1646];
                            middle <= data2[1646:1646];
                            right <= data3[1646:1646];
                        end
                    1647:
                        begin
                        left <= data1[1647:1647];
                            middle <= data2[1647:1647];
                            right <= data3[1647:1647];
                        end
                    1648:
                        begin
                        left <= data1[1648:1648];
                            middle <= data2[1648:1648];
                            right <= data3[1648:1648];
                        end
                    1649:
                        begin
                        left <= data1[1649:1649];
                            middle <= data2[1649:1649];
                            right <= data3[1649:1649];
                        end
                    1650:
                        begin
                        left <= data1[1650:1650];
                            middle <= data2[1650:1650];
                            right <= data3[1650:1650];
                        end
                    1651:
                        begin
                        left <= data1[1651:1651];
                            middle <= data2[1651:1651];
                            right <= data3[1651:1651];
                        end
                    1652:
                        begin
                        left <= data1[1652:1652];
                            middle <= data2[1652:1652];
                            right <= data3[1652:1652];
                        end
                    1653:
                        begin
                        left <= data1[1653:1653];
                            middle <= data2[1653:1653];
                            right <= data3[1653:1653];
                        end
                    1654:
                        begin
                        left <= data1[1654:1654];
                            middle <= data2[1654:1654];
                            right <= data3[1654:1654];
                        end
                    1655:
                        begin
                        left <= data1[1655:1655];
                            middle <= data2[1655:1655];
                            right <= data3[1655:1655];
                        end
                    1656:
                        begin
                        left <= data1[1656:1656];
                            middle <= data2[1656:1656];
                            right <= data3[1656:1656];
                        end
                    1657:
                        begin
                        left <= data1[1657:1657];
                            middle <= data2[1657:1657];
                            right <= data3[1657:1657];
                        end
                    1658:
                        begin
                        left <= data1[1658:1658];
                            middle <= data2[1658:1658];
                            right <= data3[1658:1658];
                        end
                    1659:
                        begin
                        left <= data1[1659:1659];
                            middle <= data2[1659:1659];
                            right <= data3[1659:1659];
                        end
                    1660:
                        begin
                        left <= data1[1660:1660];
                            middle <= data2[1660:1660];
                            right <= data3[1660:1660];
                        end
                    1661:
                        begin
                        left <= data1[1661:1661];
                            middle <= data2[1661:1661];
                            right <= data3[1661:1661];
                        end
                    1662:
                        begin
                        left <= data1[1662:1662];
                            middle <= data2[1662:1662];
                            right <= data3[1662:1662];
                        end
                    1663:
                        begin
                        left <= data1[1663:1663];
                            middle <= data2[1663:1663];
                            right <= data3[1663:1663];
                        end
                    1664:
                        begin
                        left <= data1[1664:1664];
                            middle <= data2[1664:1664];
                            right <= data3[1664:1664];
                        end
                    1665:
                        begin
                        left <= data1[1665:1665];
                            middle <= data2[1665:1665];
                            right <= data3[1665:1665];
                        end
                    1666:
                        begin
                        left <= data1[1666:1666];
                            middle <= data2[1666:1666];
                            right <= data3[1666:1666];
                        end
                    1667:
                        begin
                        left <= data1[1667:1667];
                            middle <= data2[1667:1667];
                            right <= data3[1667:1667];
                        end
                    1668:
                        begin
                        left <= data1[1668:1668];
                            middle <= data2[1668:1668];
                            right <= data3[1668:1668];
                        end
                    1669:
                        begin
                        left <= data1[1669:1669];
                            middle <= data2[1669:1669];
                            right <= data3[1669:1669];
                        end
                    1670:
                        begin
                        left <= data1[1670:1670];
                            middle <= data2[1670:1670];
                            right <= data3[1670:1670];
                        end
                    1671:
                        begin
                        left <= data1[1671:1671];
                            middle <= data2[1671:1671];
                            right <= data3[1671:1671];
                        end
                    1672:
                        begin
                        left <= data1[1672:1672];
                            middle <= data2[1672:1672];
                            right <= data3[1672:1672];
                        end
                    1673:
                        begin
                        left <= data1[1673:1673];
                            middle <= data2[1673:1673];
                            right <= data3[1673:1673];
                        end
                    1674:
                        begin
                        left <= data1[1674:1674];
                            middle <= data2[1674:1674];
                            right <= data3[1674:1674];
                        end
                    1675:
                        begin
                        left <= data1[1675:1675];
                            middle <= data2[1675:1675];
                            right <= data3[1675:1675];
                        end
                    1676:
                        begin
                        left <= data1[1676:1676];
                            middle <= data2[1676:1676];
                            right <= data3[1676:1676];
                        end
                    1677:
                        begin
                        left <= data1[1677:1677];
                            middle <= data2[1677:1677];
                            right <= data3[1677:1677];
                        end
                    1678:
                        begin
                        left <= data1[1678:1678];
                            middle <= data2[1678:1678];
                            right <= data3[1678:1678];
                        end
                    1679:
                        begin
                        left <= data1[1679:1679];
                            middle <= data2[1679:1679];
                            right <= data3[1679:1679];
                        end
                    1680:
                        begin
                        left <= data1[1680:1680];
                            middle <= data2[1680:1680];
                            right <= data3[1680:1680];
                        end
                    1681:
                        begin
                        left <= data1[1681:1681];
                            middle <= data2[1681:1681];
                            right <= data3[1681:1681];
                        end
                    1682:
                        begin
                        left <= data1[1682:1682];
                            middle <= data2[1682:1682];
                            right <= data3[1682:1682];
                        end
                    1683:
                        begin
                        left <= data1[1683:1683];
                            middle <= data2[1683:1683];
                            right <= data3[1683:1683];
                        end
                    1684:
                        begin
                        left <= data1[1684:1684];
                            middle <= data2[1684:1684];
                            right <= data3[1684:1684];
                        end
                    1685:
                        begin
                        left <= data1[1685:1685];
                            middle <= data2[1685:1685];
                            right <= data3[1685:1685];
                        end
                    1686:
                        begin
                        left <= data1[1686:1686];
                            middle <= data2[1686:1686];
                            right <= data3[1686:1686];
                        end
                    1687:
                        begin
                        left <= data1[1687:1687];
                            middle <= data2[1687:1687];
                            right <= data3[1687:1687];
                        end
                    1688:
                        begin
                        left <= data1[1688:1688];
                            middle <= data2[1688:1688];
                            right <= data3[1688:1688];
                        end
                    1689:
                        begin
                        left <= data1[1689:1689];
                            middle <= data2[1689:1689];
                            right <= data3[1689:1689];
                        end
                    1690:
                        begin
                        left <= data1[1690:1690];
                            middle <= data2[1690:1690];
                            right <= data3[1690:1690];
                        end
                    1691:
                        begin
                        left <= data1[1691:1691];
                            middle <= data2[1691:1691];
                            right <= data3[1691:1691];
                        end
                    1692:
                        begin
                        left <= data1[1692:1692];
                            middle <= data2[1692:1692];
                            right <= data3[1692:1692];
                        end
                    1693:
                        begin
                        left <= data1[1693:1693];
                            middle <= data2[1693:1693];
                            right <= data3[1693:1693];
                        end
                    1694:
                        begin
                        left <= data1[1694:1694];
                            middle <= data2[1694:1694];
                            right <= data3[1694:1694];
                        end
                    1695:
                        begin
                        left <= data1[1695:1695];
                            middle <= data2[1695:1695];
                            right <= data3[1695:1695];
                        end
                    1696:
                        begin
                        left <= data1[1696:1696];
                            middle <= data2[1696:1696];
                            right <= data3[1696:1696];
                        end
                    1697:
                        begin
                        left <= data1[1697:1697];
                            middle <= data2[1697:1697];
                            right <= data3[1697:1697];
                        end
                    1698:
                        begin
                        left <= data1[1698:1698];
                            middle <= data2[1698:1698];
                            right <= data3[1698:1698];
                        end
                    1699:
                        begin
                        left <= data1[1699:1699];
                            middle <= data2[1699:1699];
                            right <= data3[1699:1699];
                        end
                    1700:
                        begin
                        left <= data1[1700:1700];
                            middle <= data2[1700:1700];
                            right <= data3[1700:1700];
                        end
                    1701:
                        begin
                        left <= data1[1701:1701];
                            middle <= data2[1701:1701];
                            right <= data3[1701:1701];
                        end
                    1702:
                        begin
                        left <= data1[1702:1702];
                            middle <= data2[1702:1702];
                            right <= data3[1702:1702];
                        end
                    1703:
                        begin
                        left <= data1[1703:1703];
                            middle <= data2[1703:1703];
                            right <= data3[1703:1703];
                        end
                    1704:
                        begin
                        left <= data1[1704:1704];
                            middle <= data2[1704:1704];
                            right <= data3[1704:1704];
                        end
                    1705:
                        begin
                        left <= data1[1705:1705];
                            middle <= data2[1705:1705];
                            right <= data3[1705:1705];
                        end
                    1706:
                        begin
                        left <= data1[1706:1706];
                            middle <= data2[1706:1706];
                            right <= data3[1706:1706];
                        end
                    1707:
                        begin
                        left <= data1[1707:1707];
                            middle <= data2[1707:1707];
                            right <= data3[1707:1707];
                        end
                    1708:
                        begin
                        left <= data1[1708:1708];
                            middle <= data2[1708:1708];
                            right <= data3[1708:1708];
                        end
                    1709:
                        begin
                        left <= data1[1709:1709];
                            middle <= data2[1709:1709];
                            right <= data3[1709:1709];
                        end
                    1710:
                        begin
                        left <= data1[1710:1710];
                            middle <= data2[1710:1710];
                            right <= data3[1710:1710];
                        end
                    1711:
                        begin
                        left <= data1[1711:1711];
                            middle <= data2[1711:1711];
                            right <= data3[1711:1711];
                        end
                    1712:
                        begin
                        left <= data1[1712:1712];
                            middle <= data2[1712:1712];
                            right <= data3[1712:1712];
                        end
                    1713:
                        begin
                        left <= data1[1713:1713];
                            middle <= data2[1713:1713];
                            right <= data3[1713:1713];
                        end
                    1714:
                        begin
                        left <= data1[1714:1714];
                            middle <= data2[1714:1714];
                            right <= data3[1714:1714];
                        end
                    1715:
                        begin
                        left <= data1[1715:1715];
                            middle <= data2[1715:1715];
                            right <= data3[1715:1715];
                        end
                    1716:
                        begin
                        left <= data1[1716:1716];
                            middle <= data2[1716:1716];
                            right <= data3[1716:1716];
                        end
                    1717:
                        begin
                        left <= data1[1717:1717];
                            middle <= data2[1717:1717];
                            right <= data3[1717:1717];
                        end
                    1718:
                        begin
                        left <= data1[1718:1718];
                            middle <= data2[1718:1718];
                            right <= data3[1718:1718];
                        end
                    1719:
                        begin
                        left <= data1[1719:1719];
                            middle <= data2[1719:1719];
                            right <= data3[1719:1719];
                        end
                    1720:
                        begin
                        left <= data1[1720:1720];
                            middle <= data2[1720:1720];
                            right <= data3[1720:1720];
                        end
                    1721:
                        begin
                        left <= data1[1721:1721];
                            middle <= data2[1721:1721];
                            right <= data3[1721:1721];
                        end
                    1722:
                        begin
                        left <= data1[1722:1722];
                            middle <= data2[1722:1722];
                            right <= data3[1722:1722];
                        end
                    1723:
                        begin
                        left <= data1[1723:1723];
                            middle <= data2[1723:1723];
                            right <= data3[1723:1723];
                        end
                    1724:
                        begin
                        left <= data1[1724:1724];
                            middle <= data2[1724:1724];
                            right <= data3[1724:1724];
                        end
                    1725:
                        begin
                        left <= data1[1725:1725];
                            middle <= data2[1725:1725];
                            right <= data3[1725:1725];
                        end
                    1726:
                        begin
                        left <= data1[1726:1726];
                            middle <= data2[1726:1726];
                            right <= data3[1726:1726];
                        end
                    1727:
                        begin
                        left <= data1[1727:1727];
                            middle <= data2[1727:1727];
                            right <= data3[1727:1727];
                        end
                    1728:
                        begin
                        left <= data1[1728:1728];
                            middle <= data2[1728:1728];
                            right <= data3[1728:1728];
                        end
                    1729:
                        begin
                        left <= data1[1729:1729];
                            middle <= data2[1729:1729];
                            right <= data3[1729:1729];
                        end
                    1730:
                        begin
                        left <= data1[1730:1730];
                            middle <= data2[1730:1730];
                            right <= data3[1730:1730];
                        end
                    1731:
                        begin
                        left <= data1[1731:1731];
                            middle <= data2[1731:1731];
                            right <= data3[1731:1731];
                        end
                    1732:
                        begin
                        left <= data1[1732:1732];
                            middle <= data2[1732:1732];
                            right <= data3[1732:1732];
                        end
                    1733:
                        begin
                        left <= data1[1733:1733];
                            middle <= data2[1733:1733];
                            right <= data3[1733:1733];
                        end
                    1734:
                        begin
                        left <= data1[1734:1734];
                            middle <= data2[1734:1734];
                            right <= data3[1734:1734];
                        end
                    1735:
                        begin
                        left <= data1[1735:1735];
                            middle <= data2[1735:1735];
                            right <= data3[1735:1735];
                        end
                    1736:
                        begin
                        left <= data1[1736:1736];
                            middle <= data2[1736:1736];
                            right <= data3[1736:1736];
                        end
                    1737:
                        begin
                        left <= data1[1737:1737];
                            middle <= data2[1737:1737];
                            right <= data3[1737:1737];
                        end
                    1738:
                        begin
                        left <= data1[1738:1738];
                            middle <= data2[1738:1738];
                            right <= data3[1738:1738];
                        end
                    1739:
                        begin
                        left <= data1[1739:1739];
                            middle <= data2[1739:1739];
                            right <= data3[1739:1739];
                        end
                    1740:
                        begin
                        left <= data1[1740:1740];
                            middle <= data2[1740:1740];
                            right <= data3[1740:1740];
                        end
                    1741:
                        begin
                        left <= data1[1741:1741];
                            middle <= data2[1741:1741];
                            right <= data3[1741:1741];
                        end
                    1742:
                        begin
                        left <= data1[1742:1742];
                            middle <= data2[1742:1742];
                            right <= data3[1742:1742];
                        end
                    1743:
                        begin
                        left <= data1[1743:1743];
                            middle <= data2[1743:1743];
                            right <= data3[1743:1743];
                        end
                    1744:
                        begin
                        left <= data1[1744:1744];
                            middle <= data2[1744:1744];
                            right <= data3[1744:1744];
                        end
                    1745:
                        begin
                        left <= data1[1745:1745];
                            middle <= data2[1745:1745];
                            right <= data3[1745:1745];
                        end
                    1746:
                        begin
                        left <= data1[1746:1746];
                            middle <= data2[1746:1746];
                            right <= data3[1746:1746];
                        end
                    1747:
                        begin
                        left <= data1[1747:1747];
                            middle <= data2[1747:1747];
                            right <= data3[1747:1747];
                        end
                    1748:
                        begin
                        left <= data1[1748:1748];
                            middle <= data2[1748:1748];
                            right <= data3[1748:1748];
                        end
                    1749:
                        begin
                        left <= data1[1749:1749];
                            middle <= data2[1749:1749];
                            right <= data3[1749:1749];
                        end
                    1750:
                        begin
                        left <= data1[1750:1750];
                            middle <= data2[1750:1750];
                            right <= data3[1750:1750];
                        end
                    1751:
                        begin
                        left <= data1[1751:1751];
                            middle <= data2[1751:1751];
                            right <= data3[1751:1751];
                        end
                    1752:
                        begin
                        left <= data1[1752:1752];
                            middle <= data2[1752:1752];
                            right <= data3[1752:1752];
                        end
                    1753:
                        begin
                        left <= data1[1753:1753];
                            middle <= data2[1753:1753];
                            right <= data3[1753:1753];
                        end
                    1754:
                        begin
                        left <= data1[1754:1754];
                            middle <= data2[1754:1754];
                            right <= data3[1754:1754];
                        end
                    1755:
                        begin
                        left <= data1[1755:1755];
                            middle <= data2[1755:1755];
                            right <= data3[1755:1755];
                        end
                    1756:
                        begin
                        left <= data1[1756:1756];
                            middle <= data2[1756:1756];
                            right <= data3[1756:1756];
                        end
                    1757:
                        begin
                        left <= data1[1757:1757];
                            middle <= data2[1757:1757];
                            right <= data3[1757:1757];
                        end
                    1758:
                        begin
                        left <= data1[1758:1758];
                            middle <= data2[1758:1758];
                            right <= data3[1758:1758];
                        end
                    1759:
                        begin
                        left <= data1[1759:1759];
                            middle <= data2[1759:1759];
                            right <= data3[1759:1759];
                        end
                    1760:
                        begin
                        left <= data1[1760:1760];
                            middle <= data2[1760:1760];
                            right <= data3[1760:1760];
                        end
                    1761:
                        begin
                        left <= data1[1761:1761];
                            middle <= data2[1761:1761];
                            right <= data3[1761:1761];
                        end
                    1762:
                        begin
                        left <= data1[1762:1762];
                            middle <= data2[1762:1762];
                            right <= data3[1762:1762];
                        end
                    1763:
                        begin
                        left <= data1[1763:1763];
                            middle <= data2[1763:1763];
                            right <= data3[1763:1763];
                        end
                    1764:
                        begin
                        left <= data1[1764:1764];
                            middle <= data2[1764:1764];
                            right <= data3[1764:1764];
                        end
                    1765:
                        begin
                        left <= data1[1765:1765];
                            middle <= data2[1765:1765];
                            right <= data3[1765:1765];
                        end
                    1766:
                        begin
                        left <= data1[1766:1766];
                            middle <= data2[1766:1766];
                            right <= data3[1766:1766];
                        end
                    1767:
                        begin
                        left <= data1[1767:1767];
                            middle <= data2[1767:1767];
                            right <= data3[1767:1767];
                        end
                    1768:
                        begin
                        left <= data1[1768:1768];
                            middle <= data2[1768:1768];
                            right <= data3[1768:1768];
                        end
                    1769:
                        begin
                        left <= data1[1769:1769];
                            middle <= data2[1769:1769];
                            right <= data3[1769:1769];
                        end
                    1770:
                        begin
                        left <= data1[1770:1770];
                            middle <= data2[1770:1770];
                            right <= data3[1770:1770];
                        end
                    1771:
                        begin
                        left <= data1[1771:1771];
                            middle <= data2[1771:1771];
                            right <= data3[1771:1771];
                        end
                    1772:
                        begin
                        left <= data1[1772:1772];
                            middle <= data2[1772:1772];
                            right <= data3[1772:1772];
                        end
                    1773:
                        begin
                        left <= data1[1773:1773];
                            middle <= data2[1773:1773];
                            right <= data3[1773:1773];
                        end
                    1774:
                        begin
                        left <= data1[1774:1774];
                            middle <= data2[1774:1774];
                            right <= data3[1774:1774];
                        end
                    1775:
                        begin
                        left <= data1[1775:1775];
                            middle <= data2[1775:1775];
                            right <= data3[1775:1775];
                        end
                    1776:
                        begin
                        left <= data1[1776:1776];
                            middle <= data2[1776:1776];
                            right <= data3[1776:1776];
                        end
                    1777:
                        begin
                        left <= data1[1777:1777];
                            middle <= data2[1777:1777];
                            right <= data3[1777:1777];
                        end
                    1778:
                        begin
                        left <= data1[1778:1778];
                            middle <= data2[1778:1778];
                            right <= data3[1778:1778];
                        end
                    1779:
                        begin
                        left <= data1[1779:1779];
                            middle <= data2[1779:1779];
                            right <= data3[1779:1779];
                        end
                    1780:
                        begin
                        left <= data1[1780:1780];
                            middle <= data2[1780:1780];
                            right <= data3[1780:1780];
                        end
                    1781:
                        begin
                        left <= data1[1781:1781];
                            middle <= data2[1781:1781];
                            right <= data3[1781:1781];
                        end
                    1782:
                        begin
                        left <= data1[1782:1782];
                            middle <= data2[1782:1782];
                            right <= data3[1782:1782];
                        end
                    1783:
                        begin
                        left <= data1[1783:1783];
                            middle <= data2[1783:1783];
                            right <= data3[1783:1783];
                        end
                    1784:
                        begin
                        left <= data1[1784:1784];
                            middle <= data2[1784:1784];
                            right <= data3[1784:1784];
                        end
                    1785:
                        begin
                        left <= data1[1785:1785];
                            middle <= data2[1785:1785];
                            right <= data3[1785:1785];
                        end
                    1786:
                        begin
                        left <= data1[1786:1786];
                            middle <= data2[1786:1786];
                            right <= data3[1786:1786];
                        end
                    1787:
                        begin
                        left <= data1[1787:1787];
                            middle <= data2[1787:1787];
                            right <= data3[1787:1787];
                        end
                    1788:
                        begin
                        left <= data1[1788:1788];
                            middle <= data2[1788:1788];
                            right <= data3[1788:1788];
                        end
                    1789:
                        begin
                        left <= data1[1789:1789];
                            middle <= data2[1789:1789];
                            right <= data3[1789:1789];
                        end
                    1790:
                        begin
                        left <= data1[1790:1790];
                            middle <= data2[1790:1790];
                            right <= data3[1790:1790];
                        end
                    1791:
                        begin
                        left <= data1[1791:1791];
                            middle <= data2[1791:1791];
                            right <= data3[1791:1791];
                        end
                    1792:
                        begin
                        left <= data1[1792:1792];
                            middle <= data2[1792:1792];
                            right <= data3[1792:1792];
                        end
                    1793:
                        begin
                        left <= data1[1793:1793];
                            middle <= data2[1793:1793];
                            right <= data3[1793:1793];
                        end
                    1794:
                        begin
                        left <= data1[1794:1794];
                            middle <= data2[1794:1794];
                            right <= data3[1794:1794];
                        end
                    1795:
                        begin
                        left <= data1[1795:1795];
                            middle <= data2[1795:1795];
                            right <= data3[1795:1795];
                        end
                    1796:
                        begin
                        left <= data1[1796:1796];
                            middle <= data2[1796:1796];
                            right <= data3[1796:1796];
                        end
                    1797:
                        begin
                        left <= data1[1797:1797];
                            middle <= data2[1797:1797];
                            right <= data3[1797:1797];
                        end
                    1798:
                        begin
                        left <= data1[1798:1798];
                            middle <= data2[1798:1798];
                            right <= data3[1798:1798];
                        end
                    1799:
                        begin
                        left <= data1[1799:1799];
                            middle <= data2[1799:1799];
                            right <= data3[1799:1799];
                        end
                    1800:
                        begin
                        left <= data1[1800:1800];
                            middle <= data2[1800:1800];
                            right <= data3[1800:1800];
                        end
                    1801:
                        begin
                        left <= data1[1801:1801];
                            middle <= data2[1801:1801];
                            right <= data3[1801:1801];
                        end
                    1802:
                        begin
                        left <= data1[1802:1802];
                            middle <= data2[1802:1802];
                            right <= data3[1802:1802];
                        end
                    1803:
                        begin
                        left <= data1[1803:1803];
                            middle <= data2[1803:1803];
                            right <= data3[1803:1803];
                        end
                    1804:
                        begin
                        left <= data1[1804:1804];
                            middle <= data2[1804:1804];
                            right <= data3[1804:1804];
                        end
                    1805:
                        begin
                        left <= data1[1805:1805];
                            middle <= data2[1805:1805];
                            right <= data3[1805:1805];
                        end
                    1806:
                        begin
                        left <= data1[1806:1806];
                            middle <= data2[1806:1806];
                            right <= data3[1806:1806];
                        end
                    1807:
                        begin
                        left <= data1[1807:1807];
                            middle <= data2[1807:1807];
                            right <= data3[1807:1807];
                        end
                    1808:
                        begin
                        left <= data1[1808:1808];
                            middle <= data2[1808:1808];
                            right <= data3[1808:1808];
                        end
                    1809:
                        begin
                        left <= data1[1809:1809];
                            middle <= data2[1809:1809];
                            right <= data3[1809:1809];
                        end
                    1810:
                        begin
                        left <= data1[1810:1810];
                            middle <= data2[1810:1810];
                            right <= data3[1810:1810];
                        end
                    1811:
                        begin
                        left <= data1[1811:1811];
                            middle <= data2[1811:1811];
                            right <= data3[1811:1811];
                        end
                    1812:
                        begin
                        left <= data1[1812:1812];
                            middle <= data2[1812:1812];
                            right <= data3[1812:1812];
                        end
                    1813:
                        begin
                        left <= data1[1813:1813];
                            middle <= data2[1813:1813];
                            right <= data3[1813:1813];
                        end
                    1814:
                        begin
                        left <= data1[1814:1814];
                            middle <= data2[1814:1814];
                            right <= data3[1814:1814];
                        end
                    1815:
                        begin
                        left <= data1[1815:1815];
                            middle <= data2[1815:1815];
                            right <= data3[1815:1815];
                        end
                    1816:
                        begin
                        left <= data1[1816:1816];
                            middle <= data2[1816:1816];
                            right <= data3[1816:1816];
                        end
                    1817:
                        begin
                        left <= data1[1817:1817];
                            middle <= data2[1817:1817];
                            right <= data3[1817:1817];
                        end
                    1818:
                        begin
                        left <= data1[1818:1818];
                            middle <= data2[1818:1818];
                            right <= data3[1818:1818];
                        end
                    1819:
                        begin
                        left <= data1[1819:1819];
                            middle <= data2[1819:1819];
                            right <= data3[1819:1819];
                        end
                    1820:
                        begin
                        left <= data1[1820:1820];
                            middle <= data2[1820:1820];
                            right <= data3[1820:1820];
                        end
                    1821:
                        begin
                        left <= data1[1821:1821];
                            middle <= data2[1821:1821];
                            right <= data3[1821:1821];
                        end
                    1822:
                        begin
                        left <= data1[1822:1822];
                            middle <= data2[1822:1822];
                            right <= data3[1822:1822];
                        end
                    1823:
                        begin
                        left <= data1[1823:1823];
                            middle <= data2[1823:1823];
                            right <= data3[1823:1823];
                        end
                    1824:
                        begin
                        left <= data1[1824:1824];
                            middle <= data2[1824:1824];
                            right <= data3[1824:1824];
                        end
                    1825:
                        begin
                        left <= data1[1825:1825];
                            middle <= data2[1825:1825];
                            right <= data3[1825:1825];
                        end
                    1826:
                        begin
                        left <= data1[1826:1826];
                            middle <= data2[1826:1826];
                            right <= data3[1826:1826];
                        end
                    1827:
                        begin
                        left <= data1[1827:1827];
                            middle <= data2[1827:1827];
                            right <= data3[1827:1827];
                        end
                    1828:
                        begin
                        left <= data1[1828:1828];
                            middle <= data2[1828:1828];
                            right <= data3[1828:1828];
                        end
                    1829:
                        begin
                        left <= data1[1829:1829];
                            middle <= data2[1829:1829];
                            right <= data3[1829:1829];
                        end
                    1830:
                        begin
                        left <= data1[1830:1830];
                            middle <= data2[1830:1830];
                            right <= data3[1830:1830];
                        end
                    1831:
                        begin
                        left <= data1[1831:1831];
                            middle <= data2[1831:1831];
                            right <= data3[1831:1831];
                        end
                    1832:
                        begin
                        left <= data1[1832:1832];
                            middle <= data2[1832:1832];
                            right <= data3[1832:1832];
                        end
                    1833:
                        begin
                        left <= data1[1833:1833];
                            middle <= data2[1833:1833];
                            right <= data3[1833:1833];
                        end
                    1834:
                        begin
                        left <= data1[1834:1834];
                            middle <= data2[1834:1834];
                            right <= data3[1834:1834];
                        end
                    1835:
                        begin
                        left <= data1[1835:1835];
                            middle <= data2[1835:1835];
                            right <= data3[1835:1835];
                        end
                    1836:
                        begin
                        left <= data1[1836:1836];
                            middle <= data2[1836:1836];
                            right <= data3[1836:1836];
                        end
                    1837:
                        begin
                        left <= data1[1837:1837];
                            middle <= data2[1837:1837];
                            right <= data3[1837:1837];
                        end
                    1838:
                        begin
                        left <= data1[1838:1838];
                            middle <= data2[1838:1838];
                            right <= data3[1838:1838];
                        end
                    1839:
                        begin
                        left <= data1[1839:1839];
                            middle <= data2[1839:1839];
                            right <= data3[1839:1839];
                        end
                    1840:
                        begin
                        left <= data1[1840:1840];
                            middle <= data2[1840:1840];
                            right <= data3[1840:1840];
                        end
                    1841:
                        begin
                        left <= data1[1841:1841];
                            middle <= data2[1841:1841];
                            right <= data3[1841:1841];
                        end
                    1842:
                        begin
                        left <= data1[1842:1842];
                            middle <= data2[1842:1842];
                            right <= data3[1842:1842];
                        end
                    1843:
                        begin
                        left <= data1[1843:1843];
                            middle <= data2[1843:1843];
                            right <= data3[1843:1843];
                        end
                    1844:
                        begin
                        left <= data1[1844:1844];
                            middle <= data2[1844:1844];
                            right <= data3[1844:1844];
                        end
                    1845:
                        begin
                        left <= data1[1845:1845];
                            middle <= data2[1845:1845];
                            right <= data3[1845:1845];
                        end
                    1846:
                        begin
                        left <= data1[1846:1846];
                            middle <= data2[1846:1846];
                            right <= data3[1846:1846];
                        end
                    1847:
                        begin
                        left <= data1[1847:1847];
                            middle <= data2[1847:1847];
                            right <= data3[1847:1847];
                        end
                    1848:
                        begin
                        left <= data1[1848:1848];
                            middle <= data2[1848:1848];
                            right <= data3[1848:1848];
                        end
                    1849:
                        begin
                        left <= data1[1849:1849];
                            middle <= data2[1849:1849];
                            right <= data3[1849:1849];
                        end
                    1850:
                        begin
                        left <= data1[1850:1850];
                            middle <= data2[1850:1850];
                            right <= data3[1850:1850];
                        end
                    1851:
                        begin
                        left <= data1[1851:1851];
                            middle <= data2[1851:1851];
                            right <= data3[1851:1851];
                        end
                    1852:
                        begin
                        left <= data1[1852:1852];
                            middle <= data2[1852:1852];
                            right <= data3[1852:1852];
                        end
                    1853:
                        begin
                        left <= data1[1853:1853];
                            middle <= data2[1853:1853];
                            right <= data3[1853:1853];
                        end
                    1854:
                        begin
                        left <= data1[1854:1854];
                            middle <= data2[1854:1854];
                            right <= data3[1854:1854];
                        end
                    1855:
                        begin
                        left <= data1[1855:1855];
                            middle <= data2[1855:1855];
                            right <= data3[1855:1855];
                        end
                    1856:
                        begin
                        left <= data1[1856:1856];
                            middle <= data2[1856:1856];
                            right <= data3[1856:1856];
                        end
                    1857:
                        begin
                        left <= data1[1857:1857];
                            middle <= data2[1857:1857];
                            right <= data3[1857:1857];
                        end
                    1858:
                        begin
                        left <= data1[1858:1858];
                            middle <= data2[1858:1858];
                            right <= data3[1858:1858];
                        end
                    1859:
                        begin
                        left <= data1[1859:1859];
                            middle <= data2[1859:1859];
                            right <= data3[1859:1859];
                        end
                    1860:
                        begin
                        left <= data1[1860:1860];
                            middle <= data2[1860:1860];
                            right <= data3[1860:1860];
                        end
                    1861:
                        begin
                        left <= data1[1861:1861];
                            middle <= data2[1861:1861];
                            right <= data3[1861:1861];
                        end
                    1862:
                        begin
                        left <= data1[1862:1862];
                            middle <= data2[1862:1862];
                            right <= data3[1862:1862];
                        end
                    1863:
                        begin
                        left <= data1[1863:1863];
                            middle <= data2[1863:1863];
                            right <= data3[1863:1863];
                        end
                    1864:
                        begin
                        left <= data1[1864:1864];
                            middle <= data2[1864:1864];
                            right <= data3[1864:1864];
                        end
                    1865:
                        begin
                        left <= data1[1865:1865];
                            middle <= data2[1865:1865];
                            right <= data3[1865:1865];
                        end
                    1866:
                        begin
                        left <= data1[1866:1866];
                            middle <= data2[1866:1866];
                            right <= data3[1866:1866];
                        end
                    1867:
                        begin
                        left <= data1[1867:1867];
                            middle <= data2[1867:1867];
                            right <= data3[1867:1867];
                        end
                    1868:
                        begin
                        left <= data1[1868:1868];
                            middle <= data2[1868:1868];
                            right <= data3[1868:1868];
                        end
                    1869:
                        begin
                        left <= data1[1869:1869];
                            middle <= data2[1869:1869];
                            right <= data3[1869:1869];
                        end
                    1870:
                        begin
                        left <= data1[1870:1870];
                            middle <= data2[1870:1870];
                            right <= data3[1870:1870];
                        end
                    1871:
                        begin
                        left <= data1[1871:1871];
                            middle <= data2[1871:1871];
                            right <= data3[1871:1871];
                        end
                    1872:
                        begin
                        left <= data1[1872:1872];
                            middle <= data2[1872:1872];
                            right <= data3[1872:1872];
                        end
                    1873:
                        begin
                        left <= data1[1873:1873];
                            middle <= data2[1873:1873];
                            right <= data3[1873:1873];
                        end
                    1874:
                        begin
                        left <= data1[1874:1874];
                            middle <= data2[1874:1874];
                            right <= data3[1874:1874];
                        end
                    1875:
                        begin
                        left <= data1[1875:1875];
                            middle <= data2[1875:1875];
                            right <= data3[1875:1875];
                        end
                    1876:
                        begin
                        left <= data1[1876:1876];
                            middle <= data2[1876:1876];
                            right <= data3[1876:1876];
                        end
                    1877:
                        begin
                        left <= data1[1877:1877];
                            middle <= data2[1877:1877];
                            right <= data3[1877:1877];
                        end
                    1878:
                        begin
                        left <= data1[1878:1878];
                            middle <= data2[1878:1878];
                            right <= data3[1878:1878];
                        end
                    1879:
                        begin
                        left <= data1[1879:1879];
                            middle <= data2[1879:1879];
                            right <= data3[1879:1879];
                        end
                    1880:
                        begin
                        left <= data1[1880:1880];
                            middle <= data2[1880:1880];
                            right <= data3[1880:1880];
                        end
                    1881:
                        begin
                        left <= data1[1881:1881];
                            middle <= data2[1881:1881];
                            right <= data3[1881:1881];
                        end
                    1882:
                        begin
                        left <= data1[1882:1882];
                            middle <= data2[1882:1882];
                            right <= data3[1882:1882];
                        end
                    1883:
                        begin
                        left <= data1[1883:1883];
                            middle <= data2[1883:1883];
                            right <= data3[1883:1883];
                        end
                    1884:
                        begin
                        left <= data1[1884:1884];
                            middle <= data2[1884:1884];
                            right <= data3[1884:1884];
                        end
                    1885:
                        begin
                        left <= data1[1885:1885];
                            middle <= data2[1885:1885];
                            right <= data3[1885:1885];
                        end
                    1886:
                        begin
                        left <= data1[1886:1886];
                            middle <= data2[1886:1886];
                            right <= data3[1886:1886];
                        end
                    1887:
                        begin
                        left <= data1[1887:1887];
                            middle <= data2[1887:1887];
                            right <= data3[1887:1887];
                        end
                    1888:
                        begin
                        left <= data1[1888:1888];
                            middle <= data2[1888:1888];
                            right <= data3[1888:1888];
                        end
                    1889:
                        begin
                        left <= data1[1889:1889];
                            middle <= data2[1889:1889];
                            right <= data3[1889:1889];
                        end
                    1890:
                        begin
                        left <= data1[1890:1890];
                            middle <= data2[1890:1890];
                            right <= data3[1890:1890];
                        end
                    1891:
                        begin
                        left <= data1[1891:1891];
                            middle <= data2[1891:1891];
                            right <= data3[1891:1891];
                        end
                    1892:
                        begin
                        left <= data1[1892:1892];
                            middle <= data2[1892:1892];
                            right <= data3[1892:1892];
                        end
                    1893:
                        begin
                        left <= data1[1893:1893];
                            middle <= data2[1893:1893];
                            right <= data3[1893:1893];
                        end
                    1894:
                        begin
                        left <= data1[1894:1894];
                            middle <= data2[1894:1894];
                            right <= data3[1894:1894];
                        end
                    1895:
                        begin
                        left <= data1[1895:1895];
                            middle <= data2[1895:1895];
                            right <= data3[1895:1895];
                        end
                    1896:
                        begin
                        left <= data1[1896:1896];
                            middle <= data2[1896:1896];
                            right <= data3[1896:1896];
                        end
                    1897:
                        begin
                        left <= data1[1897:1897];
                            middle <= data2[1897:1897];
                            right <= data3[1897:1897];
                        end
                    1898:
                        begin
                        left <= data1[1898:1898];
                            middle <= data2[1898:1898];
                            right <= data3[1898:1898];
                        end
                    1899:
                        begin
                        left <= data1[1899:1899];
                            middle <= data2[1899:1899];
                            right <= data3[1899:1899];
                        end
                    1900:
                        begin
                        left <= data1[1900:1900];
                            middle <= data2[1900:1900];
                            right <= data3[1900:1900];
                        end
                    1901:
                        begin
                        left <= data1[1901:1901];
                            middle <= data2[1901:1901];
                            right <= data3[1901:1901];
                        end
                    1902:
                        begin
                        left <= data1[1902:1902];
                            middle <= data2[1902:1902];
                            right <= data3[1902:1902];
                        end
                    1903:
                        begin
                        left <= data1[1903:1903];
                            middle <= data2[1903:1903];
                            right <= data3[1903:1903];
                        end
                    1904:
                        begin
                        left <= data1[1904:1904];
                            middle <= data2[1904:1904];
                            right <= data3[1904:1904];
                        end
                    1905:
                        begin
                        left <= data1[1905:1905];
                            middle <= data2[1905:1905];
                            right <= data3[1905:1905];
                        end
                    1906:
                        begin
                        left <= data1[1906:1906];
                            middle <= data2[1906:1906];
                            right <= data3[1906:1906];
                        end
                    1907:
                        begin
                        left <= data1[1907:1907];
                            middle <= data2[1907:1907];
                            right <= data3[1907:1907];
                        end
                    1908:
                        begin
                        left <= data1[1908:1908];
                            middle <= data2[1908:1908];
                            right <= data3[1908:1908];
                        end
                    1909:
                        begin
                        left <= data1[1909:1909];
                            middle <= data2[1909:1909];
                            right <= data3[1909:1909];
                        end
                    1910:
                        begin
                        left <= data1[1910:1910];
                            middle <= data2[1910:1910];
                            right <= data3[1910:1910];
                        end
                    1911:
                        begin
                        left <= data1[1911:1911];
                            middle <= data2[1911:1911];
                            right <= data3[1911:1911];
                        end
                    1912:
                        begin
                        left <= data1[1912:1912];
                            middle <= data2[1912:1912];
                            right <= data3[1912:1912];
                        end
                    1913:
                        begin
                        left <= data1[1913:1913];
                            middle <= data2[1913:1913];
                            right <= data3[1913:1913];
                        end
                    1914:
                        begin
                        left <= data1[1914:1914];
                            middle <= data2[1914:1914];
                            right <= data3[1914:1914];
                        end
                    1915:
                        begin
                        left <= data1[1915:1915];
                            middle <= data2[1915:1915];
                            right <= data3[1915:1915];
                        end
                    1916:
                        begin
                        left <= data1[1916:1916];
                            middle <= data2[1916:1916];
                            right <= data3[1916:1916];
                        end
                    1917:
                        begin
                        left <= data1[1917:1917];
                            middle <= data2[1917:1917];
                            right <= data3[1917:1917];
                        end
                    1918:
                        begin
                        left <= data1[1918:1918];
                            middle <= data2[1918:1918];
                            right <= data3[1918:1918];
                        end
                    1919:
                        begin
                        left <= data1[1919:1919];
                            middle <= data2[1919:1919];
                            right <= data3[1919:1919];
                        end
                    1920:
                        begin
                        left <= data1[1920:1920];
                            middle <= data2[1920:1920];
                            right <= data3[1920:1920];
                        end
                    1921:
                        begin
                        left <= data1[1921:1921];
                            middle <= data2[1921:1921];
                            right <= data3[1921:1921];
                        end
                    1922:
                        begin
                        left <= data1[1922:1922];
                            middle <= data2[1922:1922];
                            right <= data3[1922:1922];
                        end
                    1923:
                        begin
                        left <= data1[1923:1923];
                            middle <= data2[1923:1923];
                            right <= data3[1923:1923];
                        end
                    1924:
                        begin
                        left <= data1[1924:1924];
                            middle <= data2[1924:1924];
                            right <= data3[1924:1924];
                        end
                    1925:
                        begin
                        left <= data1[1925:1925];
                            middle <= data2[1925:1925];
                            right <= data3[1925:1925];
                        end
                    1926:
                        begin
                        left <= data1[1926:1926];
                            middle <= data2[1926:1926];
                            right <= data3[1926:1926];
                        end
                    1927:
                        begin
                        left <= data1[1927:1927];
                            middle <= data2[1927:1927];
                            right <= data3[1927:1927];
                        end
                    1928:
                        begin
                        left <= data1[1928:1928];
                            middle <= data2[1928:1928];
                            right <= data3[1928:1928];
                        end
                    1929:
                        begin
                        left <= data1[1929:1929];
                            middle <= data2[1929:1929];
                            right <= data3[1929:1929];
                        end
                    1930:
                        begin
                        left <= data1[1930:1930];
                            middle <= data2[1930:1930];
                            right <= data3[1930:1930];
                        end
                    1931:
                        begin
                        left <= data1[1931:1931];
                            middle <= data2[1931:1931];
                            right <= data3[1931:1931];
                        end
                    1932:
                        begin
                        left <= data1[1932:1932];
                            middle <= data2[1932:1932];
                            right <= data3[1932:1932];
                        end
                    1933:
                        begin
                        left <= data1[1933:1933];
                            middle <= data2[1933:1933];
                            right <= data3[1933:1933];
                        end
                    1934:
                        begin
                        left <= data1[1934:1934];
                            middle <= data2[1934:1934];
                            right <= data3[1934:1934];
                        end
                    1935:
                        begin
                        left <= data1[1935:1935];
                            middle <= data2[1935:1935];
                            right <= data3[1935:1935];
                        end
                    1936:
                        begin
                        left <= data1[1936:1936];
                            middle <= data2[1936:1936];
                            right <= data3[1936:1936];
                        end
                    1937:
                        begin
                        left <= data1[1937:1937];
                            middle <= data2[1937:1937];
                            right <= data3[1937:1937];
                        end
                    1938:
                        begin
                        left <= data1[1938:1938];
                            middle <= data2[1938:1938];
                            right <= data3[1938:1938];
                        end
                    1939:
                        begin
                        left <= data1[1939:1939];
                            middle <= data2[1939:1939];
                            right <= data3[1939:1939];
                        end
                    1940:
                        begin
                        left <= data1[1940:1940];
                            middle <= data2[1940:1940];
                            right <= data3[1940:1940];
                        end
                    1941:
                        begin
                        left <= data1[1941:1941];
                            middle <= data2[1941:1941];
                            right <= data3[1941:1941];
                        end
                    1942:
                        begin
                        left <= data1[1942:1942];
                            middle <= data2[1942:1942];
                            right <= data3[1942:1942];
                        end
                    1943:
                        begin
                        left <= data1[1943:1943];
                            middle <= data2[1943:1943];
                            right <= data3[1943:1943];
                        end
                    1944:
                        begin
                        left <= data1[1944:1944];
                            middle <= data2[1944:1944];
                            right <= data3[1944:1944];
                        end
                    1945:
                        begin
                        left <= data1[1945:1945];
                            middle <= data2[1945:1945];
                            right <= data3[1945:1945];
                        end
                    1946:
                        begin
                        left <= data1[1946:1946];
                            middle <= data2[1946:1946];
                            right <= data3[1946:1946];
                        end
                    1947:
                        begin
                        left <= data1[1947:1947];
                            middle <= data2[1947:1947];
                            right <= data3[1947:1947];
                        end
                    1948:
                        begin
                        left <= data1[1948:1948];
                            middle <= data2[1948:1948];
                            right <= data3[1948:1948];
                        end
                    1949:
                        begin
                        left <= data1[1949:1949];
                            middle <= data2[1949:1949];
                            right <= data3[1949:1949];
                        end
                    1950:
                        begin
                        left <= data1[1950:1950];
                            middle <= data2[1950:1950];
                            right <= data3[1950:1950];
                        end
                    1951:
                        begin
                        left <= data1[1951:1951];
                            middle <= data2[1951:1951];
                            right <= data3[1951:1951];
                        end
                    1952:
                        begin
                        left <= data1[1952:1952];
                            middle <= data2[1952:1952];
                            right <= data3[1952:1952];
                        end
                    1953:
                        begin
                        left <= data1[1953:1953];
                            middle <= data2[1953:1953];
                            right <= data3[1953:1953];
                        end
                    1954:
                        begin
                        left <= data1[1954:1954];
                            middle <= data2[1954:1954];
                            right <= data3[1954:1954];
                        end
                    1955:
                        begin
                        left <= data1[1955:1955];
                            middle <= data2[1955:1955];
                            right <= data3[1955:1955];
                        end
                    1956:
                        begin
                        left <= data1[1956:1956];
                            middle <= data2[1956:1956];
                            right <= data3[1956:1956];
                        end
                    1957:
                        begin
                        left <= data1[1957:1957];
                            middle <= data2[1957:1957];
                            right <= data3[1957:1957];
                        end
                    1958:
                        begin
                        left <= data1[1958:1958];
                            middle <= data2[1958:1958];
                            right <= data3[1958:1958];
                        end
                    1959:
                        begin
                        left <= data1[1959:1959];
                            middle <= data2[1959:1959];
                            right <= data3[1959:1959];
                        end
                    1960:
                        begin
                        left <= data1[1960:1960];
                            middle <= data2[1960:1960];
                            right <= data3[1960:1960];
                        end
                    1961:
                        begin
                        left <= data1[1961:1961];
                            middle <= data2[1961:1961];
                            right <= data3[1961:1961];
                        end
                    1962:
                        begin
                        left <= data1[1962:1962];
                            middle <= data2[1962:1962];
                            right <= data3[1962:1962];
                        end
                    1963:
                        begin
                        left <= data1[1963:1963];
                            middle <= data2[1963:1963];
                            right <= data3[1963:1963];
                        end
                    1964:
                        begin
                        left <= data1[1964:1964];
                            middle <= data2[1964:1964];
                            right <= data3[1964:1964];
                        end
                    1965:
                        begin
                        left <= data1[1965:1965];
                            middle <= data2[1965:1965];
                            right <= data3[1965:1965];
                        end
                    1966:
                        begin
                        left <= data1[1966:1966];
                            middle <= data2[1966:1966];
                            right <= data3[1966:1966];
                        end
                    1967:
                        begin
                        left <= data1[1967:1967];
                            middle <= data2[1967:1967];
                            right <= data3[1967:1967];
                        end
                    1968:
                        begin
                        left <= data1[1968:1968];
                            middle <= data2[1968:1968];
                            right <= data3[1968:1968];
                        end
                    1969:
                        begin
                        left <= data1[1969:1969];
                            middle <= data2[1969:1969];
                            right <= data3[1969:1969];
                        end
                    1970:
                        begin
                        left <= data1[1970:1970];
                            middle <= data2[1970:1970];
                            right <= data3[1970:1970];
                        end
                    1971:
                        begin
                        left <= data1[1971:1971];
                            middle <= data2[1971:1971];
                            right <= data3[1971:1971];
                        end
                    1972:
                        begin
                        left <= data1[1972:1972];
                            middle <= data2[1972:1972];
                            right <= data3[1972:1972];
                        end
                    1973:
                        begin
                        left <= data1[1973:1973];
                            middle <= data2[1973:1973];
                            right <= data3[1973:1973];
                        end
                    1974:
                        begin
                        left <= data1[1974:1974];
                            middle <= data2[1974:1974];
                            right <= data3[1974:1974];
                        end
                    1975:
                        begin
                        left <= data1[1975:1975];
                            middle <= data2[1975:1975];
                            right <= data3[1975:1975];
                        end
                    1976:
                        begin
                        left <= data1[1976:1976];
                            middle <= data2[1976:1976];
                            right <= data3[1976:1976];
                        end
                    1977:
                        begin
                        left <= data1[1977:1977];
                            middle <= data2[1977:1977];
                            right <= data3[1977:1977];
                        end
                    1978:
                        begin
                        left <= data1[1978:1978];
                            middle <= data2[1978:1978];
                            right <= data3[1978:1978];
                        end
                    1979:
                        begin
                        left <= data1[1979:1979];
                            middle <= data2[1979:1979];
                            right <= data3[1979:1979];
                        end
                    1980:
                        begin
                        left <= data1[1980:1980];
                            middle <= data2[1980:1980];
                            right <= data3[1980:1980];
                        end
                    1981:
                        begin
                        left <= data1[1981:1981];
                            middle <= data2[1981:1981];
                            right <= data3[1981:1981];
                        end
                    1982:
                        begin
                        left <= data1[1982:1982];
                            middle <= data2[1982:1982];
                            right <= data3[1982:1982];
                        end
                    1983:
                        begin
                        left <= data1[1983:1983];
                            middle <= data2[1983:1983];
                            right <= data3[1983:1983];
                        end
                    1984:
                        begin
                        left <= data1[1984:1984];
                            middle <= data2[1984:1984];
                            right <= data3[1984:1984];
                        end
                    1985:
                        begin
                        left <= data1[1985:1985];
                            middle <= data2[1985:1985];
                            right <= data3[1985:1985];
                        end
                    1986:
                        begin
                        left <= data1[1986:1986];
                            middle <= data2[1986:1986];
                            right <= data3[1986:1986];
                        end
                    1987:
                        begin
                        left <= data1[1987:1987];
                            middle <= data2[1987:1987];
                            right <= data3[1987:1987];
                        end
                    1988:
                        begin
                        left <= data1[1988:1988];
                            middle <= data2[1988:1988];
                            right <= data3[1988:1988];
                        end
                    1989:
                        begin
                        left <= data1[1989:1989];
                            middle <= data2[1989:1989];
                            right <= data3[1989:1989];
                        end
                    1990:
                        begin
                        left <= data1[1990:1990];
                            middle <= data2[1990:1990];
                            right <= data3[1990:1990];
                        end
                    1991:
                        begin
                        left <= data1[1991:1991];
                            middle <= data2[1991:1991];
                            right <= data3[1991:1991];
                        end
                    1992:
                        begin
                        left <= data1[1992:1992];
                            middle <= data2[1992:1992];
                            right <= data3[1992:1992];
                        end
                    1993:
                        begin
                        left <= data1[1993:1993];
                            middle <= data2[1993:1993];
                            right <= data3[1993:1993];
                        end
                    1994:
                        begin
                        left <= data1[1994:1994];
                            middle <= data2[1994:1994];
                            right <= data3[1994:1994];
                        end
                    1995:
                        begin
                        left <= data1[1995:1995];
                            middle <= data2[1995:1995];
                            right <= data3[1995:1995];
                        end
                    1996:
                        begin
                        left <= data1[1996:1996];
                            middle <= data2[1996:1996];
                            right <= data3[1996:1996];
                        end
                    1997:
                        begin
                        left <= data1[1997:1997];
                            middle <= data2[1997:1997];
                            right <= data3[1997:1997];
                        end
                    1998:
                        begin
                        left <= data1[1998:1998];
                            middle <= data2[1998:1998];
                            right <= data3[1998:1998];
                        end
                    1999:
                        begin
                        left <= data1[1999:1999];
                            middle <= data2[1999:1999];
                            right <= data3[1999:1999];
                        end
                    2000:
                        begin
                        left <= data1[2000:2000];
                            middle <= data2[2000:2000];
                            right <= data3[2000:2000];
                        end
                    2001:
                        begin
                        left <= data1[2001:2001];
                            middle <= data2[2001:2001];
                            right <= data3[2001:2001];
                        end
                    2002:
                        begin
                        left <= data1[2002:2002];
                            middle <= data2[2002:2002];
                            right <= data3[2002:2002];
                        end
                    2003:
                        begin
                        left <= data1[2003:2003];
                            middle <= data2[2003:2003];
                            right <= data3[2003:2003];
                        end
                    2004:
                        begin
                        left <= data1[2004:2004];
                            middle <= data2[2004:2004];
                            right <= data3[2004:2004];
                        end
                    2005:
                        begin
                        left <= data1[2005:2005];
                            middle <= data2[2005:2005];
                            right <= data3[2005:2005];
                        end
                    2006:
                        begin
                        left <= data1[2006:2006];
                            middle <= data2[2006:2006];
                            right <= data3[2006:2006];
                        end
                    2007:
                        begin
                        left <= data1[2007:2007];
                            middle <= data2[2007:2007];
                            right <= data3[2007:2007];
                        end
                    2008:
                        begin
                        left <= data1[2008:2008];
                            middle <= data2[2008:2008];
                            right <= data3[2008:2008];
                        end
                    2009:
                        begin
                        left <= data1[2009:2009];
                            middle <= data2[2009:2009];
                            right <= data3[2009:2009];
                        end
                    2010:
                        begin
                        left <= data1[2010:2010];
                            middle <= data2[2010:2010];
                            right <= data3[2010:2010];
                        end
                    2011:
                        begin
                        left <= data1[2011:2011];
                            middle <= data2[2011:2011];
                            right <= data3[2011:2011];
                        end
                    2012:
                        begin
                        left <= data1[2012:2012];
                            middle <= data2[2012:2012];
                            right <= data3[2012:2012];
                        end
                    2013:
                        begin
                        left <= data1[2013:2013];
                            middle <= data2[2013:2013];
                            right <= data3[2013:2013];
                        end
                    2014:
                        begin
                        left <= data1[2014:2014];
                            middle <= data2[2014:2014];
                            right <= data3[2014:2014];
                        end
                    2015:
                        begin
                        left <= data1[2015:2015];
                            middle <= data2[2015:2015];
                            right <= data3[2015:2015];
                        end
                    2016:
                        begin
                        left <= data1[2016:2016];
                            middle <= data2[2016:2016];
                            right <= data3[2016:2016];
                        end
                    2017:
                        begin
                        left <= data1[2017:2017];
                            middle <= data2[2017:2017];
                            right <= data3[2017:2017];
                        end
                    2018:
                        begin
                        left <= data1[2018:2018];
                            middle <= data2[2018:2018];
                            right <= data3[2018:2018];
                        end
                    2019:
                        begin
                        left <= data1[2019:2019];
                            middle <= data2[2019:2019];
                            right <= data3[2019:2019];
                        end
                    2020:
                        begin
                        left <= data1[2020:2020];
                            middle <= data2[2020:2020];
                            right <= data3[2020:2020];
                        end
                    2021:
                        begin
                        left <= data1[2021:2021];
                            middle <= data2[2021:2021];
                            right <= data3[2021:2021];
                        end
                    2022:
                        begin
                        left <= data1[2022:2022];
                            middle <= data2[2022:2022];
                            right <= data3[2022:2022];
                        end
                    2023:
                        begin
                        left <= data1[2023:2023];
                            middle <= data2[2023:2023];
                            right <= data3[2023:2023];
                        end
                    2024:
                        begin
                        left <= data1[2024:2024];
                            middle <= data2[2024:2024];
                            right <= data3[2024:2024];
                        end
                    2025:
                        begin
                        left <= data1[2025:2025];
                            middle <= data2[2025:2025];
                            right <= data3[2025:2025];
                        end
                    2026:
                        begin
                        left <= data1[2026:2026];
                            middle <= data2[2026:2026];
                            right <= data3[2026:2026];
                        end
                    2027:
                        begin
                        left <= data1[2027:2027];
                            middle <= data2[2027:2027];
                            right <= data3[2027:2027];
                        end
                    2028:
                        begin
                        left <= data1[2028:2028];
                            middle <= data2[2028:2028];
                            right <= data3[2028:2028];
                        end
                    2029:
                        begin
                        left <= data1[2029:2029];
                            middle <= data2[2029:2029];
                            right <= data3[2029:2029];
                        end
                    2030:
                        begin
                        left <= data1[2030:2030];
                            middle <= data2[2030:2030];
                            right <= data3[2030:2030];
                        end
                    2031:
                        begin
                        left <= data1[2031:2031];
                            middle <= data2[2031:2031];
                            right <= data3[2031:2031];
                        end
                    2032:
                        begin
                        left <= data1[2032:2032];
                            middle <= data2[2032:2032];
                            right <= data3[2032:2032];
                        end
                    2033:
                        begin
                        left <= data1[2033:2033];
                            middle <= data2[2033:2033];
                            right <= data3[2033:2033];
                        end
                    2034:
                        begin
                        left <= data1[2034:2034];
                            middle <= data2[2034:2034];
                            right <= data3[2034:2034];
                        end
                    2035:
                        begin
                        left <= data1[2035:2035];
                            middle <= data2[2035:2035];
                            right <= data3[2035:2035];
                        end
                    2036:
                        begin
                        left <= data1[2036:2036];
                            middle <= data2[2036:2036];
                            right <= data3[2036:2036];
                        end
                    2037:
                        begin
                        left <= data1[2037:2037];
                            middle <= data2[2037:2037];
                            right <= data3[2037:2037];
                        end
                    2038:
                        begin
                        left <= data1[2038:2038];
                            middle <= data2[2038:2038];
                            right <= data3[2038:2038];
                        end
                    2039:
                        begin
                        left <= data1[2039:2039];
                            middle <= data2[2039:2039];
                            right <= data3[2039:2039];
                        end
                    2040:
                        begin
                        left <= data1[2040:2040];
                            middle <= data2[2040:2040];
                            right <= data3[2040:2040];
                        end
                    2041:
                        begin
                        left <= data1[2041:2041];
                            middle <= data2[2041:2041];
                            right <= data3[2041:2041];
                        end
                    2042:
                        begin
                        left <= data1[2042:2042];
                            middle <= data2[2042:2042];
                            right <= data3[2042:2042];
                        end
                    2043:
                        begin
                        left <= data1[2043:2043];
                            middle <= data2[2043:2043];
                            right <= data3[2043:2043];
                        end
                    2044:
                        begin
                        left <= data1[2044:2044];
                            middle <= data2[2044:2044];
                            right <= data3[2044:2044];
                        end
                    2045:
                        begin
                        left <= data1[2045:2045];
                            middle <= data2[2045:2045];
                            right <= data3[2045:2045];
                        end
                    2046:
                        begin
                        left <= data1[2046:2046];
                            middle <= data2[2046:2046];
                            right <= data3[2046:2046];
                        end
                    2047:
                        begin
                        left <= data1[2047:2047];
                            middle <= data2[2047:2047];
                            right <= data3[2047:2047];
                        end
                endcase

				show0[6:0] = show1[6:0];
				show1[6:0] = show2[6:0];
				show2[6:0] = show3[6:0];
				show3[6:0] = show4[6:0];
				show4[6:0] = show5[6:0];
				show5[6:0] = {~middle, 2'b11, ~right, 2'b11, ~left};
				end
			end
		end
	end

	generator_1000hz(c, clk);
	counter_scan(clk, scan_cnt);
	selector_digit(scan_cnt, SEGNum);
	selector_seg(scan_cnt, show0, show1, show2, show3, show4, show5, L);

endmodule